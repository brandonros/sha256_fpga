// synchronous circuit fpga_test::Sha256Core
module top(input wire [1:0] clock_reset, input wire [512:0] i, output wire [0:0] o);
    wire [1153:0] od;
    wire [1152:0] d;
    wire [1152:0] q;
    assign o = od[0];
    top_state c0 (.clock_reset(clock_reset),.i(d[640:0]),.o(q[640:0]));
    top_w c1 (.clock_reset(clock_reset),.i(d[1152:641]),.o(q[1152:641]));
    assign od = kernel_kernel(clock_reset, i, q);
    assign d = od[1153:1];
    function [1153:0] kernel_kernel(input reg [1:0] arg_0, input reg [512:0] arg_1, input reg [1152:0] arg_2);
        reg [0:0] r0;
        reg [512:0] r1;
        reg [511:0] r2;
        reg [31:0] r3;
        reg [1152:0] r4;
        reg [511:0] r5;
        reg [31:0] r6;
        reg [1152:0] r7;
        reg [511:0] r8;
        reg [31:0] r9;
        reg [1152:0] r10;
        reg [511:0] r11;
        reg [31:0] r12;
        reg [1152:0] r13;
        reg [511:0] r14;
        reg [31:0] r15;
        reg [1152:0] r16;
        reg [511:0] r17;
        reg [31:0] r18;
        reg [1152:0] r19;
        reg [511:0] r20;
        reg [31:0] r21;
        reg [1152:0] r22;
        reg [511:0] r23;
        reg [31:0] r24;
        reg [1152:0] r25;
        reg [511:0] r26;
        reg [31:0] r27;
        reg [1152:0] r28;
        reg [511:0] r29;
        reg [31:0] r30;
        reg [1152:0] r31;
        reg [511:0] r32;
        reg [31:0] r33;
        reg [1152:0] r34;
        reg [511:0] r35;
        reg [31:0] r36;
        reg [1152:0] r37;
        reg [511:0] r38;
        reg [31:0] r39;
        reg [1152:0] r40;
        reg [511:0] r41;
        reg [31:0] r42;
        reg [1152:0] r43;
        reg [511:0] r44;
        reg [31:0] r45;
        reg [1152:0] r46;
        reg [511:0] r47;
        reg [31:0] r48;
        reg [1152:0] r49;
        reg [640:0] r50;
        reg [1152:0] r51;
        reg [0:0] r52;
        reg [0:0] r53;
        reg [640:0] r54;
        reg [127:0] r55;
        reg [640:0] r56;
        reg [1152:0] r57;
        reg [0:0] r58;
        reg [511:0] r59;
        reg [31:0] r60;
        reg [1152:0] r61;
        reg [511:0] r62;
        reg [31:0] r63;
        reg [1152:0] r64;
        reg [511:0] r65;
        reg [31:0] r66;
        reg [1152:0] r67;
        reg [511:0] r68;
        reg [31:0] r69;
        reg [1152:0] r70;
        reg [511:0] r71;
        reg [31:0] r72;
        reg [1152:0] r73;
        reg [511:0] r74;
        reg [31:0] r75;
        reg [1152:0] r76;
        reg [511:0] r77;
        reg [31:0] r78;
        reg [1152:0] r79;
        reg [511:0] r80;
        reg [31:0] r81;
        reg [1152:0] r82;
        reg [511:0] r83;
        reg [31:0] r84;
        reg [1152:0] r85;
        reg [511:0] r86;
        reg [31:0] r87;
        reg [1152:0] r88;
        reg [511:0] r89;
        reg [31:0] r90;
        reg [1152:0] r91;
        reg [511:0] r92;
        reg [31:0] r93;
        reg [1152:0] r94;
        reg [511:0] r95;
        reg [31:0] r96;
        reg [1152:0] r97;
        reg [511:0] r98;
        reg [31:0] r99;
        reg [1152:0] r100;
        reg [511:0] r101;
        reg [31:0] r102;
        reg [1152:0] r103;
        reg [640:0] r104;
        reg [127:0] r105;
        reg [511:0] r106;
        reg [31:0] r107;
        reg [511:0] r108;
        reg [31:0] r109;
        reg [511:0] r110;
        reg [31:0] r111;
        reg [511:0] r112;
        reg [31:0] r113;
        reg [31:0] r119;
        reg [0:0] r120;
        reg [31:0] r125;
        reg [31:0] r127;
        reg [31:0] r128;
        reg [31:0] r133;
        reg [31:0] r135;
        reg [31:0] r136;
        reg [31:0] r138;
        reg [31:0] r139;
        reg [31:0] r140;
        reg [31:0] r142;
        reg [31:0] r147;
        reg [31:0] r149;
        reg [31:0] r150;
        reg [31:0] r155;
        reg [31:0] r157;
        reg [31:0] r158;
        reg [31:0] r160;
        reg [31:0] r161;
        reg [31:0] r162;
        reg [31:0] r164;
        reg [31:0] r165;
        reg [1152:0] r167;
        reg [511:0] r168;
        reg [31:0] r169;
        reg [1152:0] r170;
        reg [511:0] r171;
        reg [31:0] r172;
        reg [1152:0] r173;
        reg [511:0] r174;
        reg [31:0] r175;
        reg [1152:0] r176;
        reg [511:0] r177;
        reg [31:0] r178;
        reg [1152:0] r179;
        reg [511:0] r180;
        reg [31:0] r181;
        reg [1152:0] r182;
        reg [511:0] r183;
        reg [31:0] r184;
        reg [1152:0] r185;
        reg [511:0] r186;
        reg [31:0] r187;
        reg [1152:0] r188;
        reg [511:0] r189;
        reg [31:0] r190;
        reg [1152:0] r191;
        reg [511:0] r192;
        reg [31:0] r193;
        reg [1152:0] r194;
        reg [511:0] r195;
        reg [31:0] r196;
        reg [1152:0] r197;
        reg [511:0] r198;
        reg [31:0] r199;
        reg [1152:0] r200;
        reg [511:0] r201;
        reg [31:0] r202;
        reg [1152:0] r203;
        reg [511:0] r204;
        reg [31:0] r205;
        reg [1152:0] r206;
        reg [511:0] r207;
        reg [31:0] r208;
        reg [1152:0] r209;
        reg [511:0] r210;
        reg [31:0] r211;
        reg [1152:0] r212;
        reg [511:0] r213;
        reg [31:0] r214;
        reg [1152:0] r215;
        reg [1152:0] r216;
        reg [0:0] r217;
        reg [0:0] r218;
        reg [63:0] r219;
        reg [0:0] r220;
        reg [511:0] r221;
        reg [31:0] r222;
        reg [0:0] r223;
        reg [511:0] r224;
        reg [31:0] r225;
        reg [0:0] r226;
        reg [511:0] r227;
        reg [31:0] r228;
        reg [0:0] r229;
        reg [511:0] r230;
        reg [31:0] r231;
        reg [0:0] r232;
        reg [511:0] r233;
        reg [31:0] r234;
        reg [0:0] r235;
        reg [511:0] r236;
        reg [31:0] r237;
        reg [0:0] r238;
        reg [511:0] r239;
        reg [31:0] r240;
        reg [0:0] r241;
        reg [511:0] r242;
        reg [31:0] r243;
        reg [0:0] r244;
        reg [511:0] r245;
        reg [31:0] r246;
        reg [0:0] r247;
        reg [511:0] r248;
        reg [31:0] r249;
        reg [0:0] r250;
        reg [511:0] r251;
        reg [31:0] r252;
        reg [0:0] r253;
        reg [511:0] r254;
        reg [31:0] r255;
        reg [0:0] r256;
        reg [511:0] r257;
        reg [31:0] r258;
        reg [0:0] r259;
        reg [511:0] r260;
        reg [31:0] r261;
        reg [0:0] r262;
        reg [511:0] r263;
        reg [31:0] r264;
        reg [511:0] r265;
        reg [31:0] r266;
        reg [31:0] r267;
        reg [31:0] r268;
        reg [31:0] r269;
        reg [31:0] r270;
        reg [31:0] r271;
        reg [31:0] r272;
        reg [31:0] r273;
        reg [31:0] r274;
        reg [31:0] r275;
        reg [31:0] r276;
        reg [31:0] r277;
        reg [31:0] r278;
        reg [31:0] r279;
        reg [31:0] r280;
        reg [31:0] r281;
        reg [511:0] r282;
        reg [31:0] r283;
        reg [31:0] r284;
        reg [640:0] r285;
        reg [31:0] r286;
        reg [31:0] r288;
        reg [31:0] r292;
        reg [31:0] r294;
        reg [31:0] r295;
        reg [31:0] r300;
        reg [31:0] r302;
        reg [31:0] r303;
        reg [31:0] r305;
        reg [31:0] r309;
        reg [31:0] r311;
        reg [31:0] r312;
        reg [640:0] r315;
        reg [31:0] r316;
        reg [640:0] r317;
        reg [31:0] r318;
        reg [640:0] r319;
        reg [31:0] r320;
        reg [31:0] r324;
        reg [31:0] r325;
        reg [31:0] r326;
        reg [31:0] r327;
        reg [640:0] r329;
        reg [31:0] r330;
        reg [31:0] r331;
        reg [31:0] r332;
        reg [640:0] r333;
        reg [127:0] r334;
        reg [31:0] r336;
        reg [63:0] r337;
        reg [0:0] r338;
        reg [13:0] r339;
        reg [27:0] r340;
        reg [13:0] r341;
        reg [13:0] r342;
        reg [127:0] r343;
        reg [31:0] r344;
        reg [31:0] r346;
        reg [31:0] r347;
        reg [640:0] r348;
        reg [31:0] r349;
        reg [31:0] r351;
        reg [31:0] r355;
        reg [31:0] r357;
        reg [31:0] r358;
        reg [31:0] r363;
        reg [31:0] r365;
        reg [31:0] r366;
        reg [31:0] r368;
        reg [31:0] r372;
        reg [31:0] r374;
        reg [31:0] r375;
        reg [640:0] r378;
        reg [31:0] r379;
        reg [640:0] r380;
        reg [31:0] r381;
        reg [640:0] r382;
        reg [31:0] r383;
        reg [31:0] r387;
        reg [31:0] r388;
        reg [31:0] r389;
        reg [31:0] r390;
        reg [31:0] r391;
        reg [31:0] r393;
        reg [640:0] r394;
        reg [31:0] r395;
        reg [1152:0] r396;
        reg [640:0] r397;
        reg [31:0] r398;
        reg [1152:0] r399;
        reg [640:0] r400;
        reg [31:0] r401;
        reg [1152:0] r402;
        reg [640:0] r403;
        reg [31:0] r404;
        reg [31:0] r405;
        reg [1152:0] r406;
        reg [640:0] r407;
        reg [31:0] r408;
        reg [1152:0] r409;
        reg [640:0] r410;
        reg [31:0] r411;
        reg [1152:0] r412;
        reg [640:0] r413;
        reg [31:0] r414;
        reg [1152:0] r415;
        reg [31:0] r416;
        reg [1152:0] r417;
        reg [127:0] r418;
        reg [127:0] r419;
        reg [1152:0] r420;
        reg [0:0] r421;
        reg [640:0] r422;
        reg [255:0] r423;
        reg [31:0] r424;
        reg [640:0] r425;
        reg [31:0] r426;
        reg [31:0] r427;
        reg [1152:0] r428;
        reg [640:0] r429;
        reg [255:0] r430;
        reg [31:0] r431;
        reg [640:0] r432;
        reg [31:0] r433;
        reg [31:0] r434;
        reg [1152:0] r435;
        reg [640:0] r436;
        reg [255:0] r437;
        reg [31:0] r438;
        reg [640:0] r439;
        reg [31:0] r440;
        reg [31:0] r441;
        reg [1152:0] r442;
        reg [640:0] r443;
        reg [255:0] r444;
        reg [31:0] r445;
        reg [640:0] r446;
        reg [31:0] r447;
        reg [31:0] r448;
        reg [1152:0] r449;
        reg [640:0] r450;
        reg [255:0] r451;
        reg [31:0] r452;
        reg [640:0] r453;
        reg [31:0] r454;
        reg [31:0] r455;
        reg [1152:0] r456;
        reg [640:0] r457;
        reg [255:0] r458;
        reg [31:0] r459;
        reg [640:0] r460;
        reg [31:0] r461;
        reg [31:0] r462;
        reg [1152:0] r463;
        reg [640:0] r464;
        reg [255:0] r465;
        reg [31:0] r466;
        reg [640:0] r467;
        reg [31:0] r468;
        reg [31:0] r469;
        reg [1152:0] r470;
        reg [640:0] r471;
        reg [255:0] r472;
        reg [31:0] r473;
        reg [640:0] r474;
        reg [31:0] r475;
        reg [31:0] r476;
        reg [1152:0] r477;
        reg [1152:0] r478;
        reg [1152:0] r479;
        reg [1152:0] r480;
        reg [640:0] r481;
        reg [1152:0] r482;
        reg [511:0] r483;
        reg [31:0] r484;
        reg [1152:0] r485;
        reg [511:0] r486;
        reg [31:0] r487;
        reg [1152:0] r488;
        reg [511:0] r489;
        reg [31:0] r490;
        reg [1152:0] r491;
        reg [511:0] r492;
        reg [31:0] r493;
        reg [1152:0] r494;
        reg [511:0] r495;
        reg [31:0] r496;
        reg [1152:0] r497;
        reg [511:0] r498;
        reg [31:0] r499;
        reg [1152:0] r500;
        reg [511:0] r501;
        reg [31:0] r502;
        reg [1152:0] r503;
        reg [511:0] r504;
        reg [31:0] r505;
        reg [1152:0] r506;
        reg [511:0] r507;
        reg [31:0] r508;
        reg [1152:0] r509;
        reg [511:0] r510;
        reg [31:0] r511;
        reg [1152:0] r512;
        reg [511:0] r513;
        reg [31:0] r514;
        reg [1152:0] r515;
        reg [511:0] r516;
        reg [31:0] r517;
        reg [1152:0] r518;
        reg [511:0] r519;
        reg [31:0] r520;
        reg [1152:0] r521;
        reg [511:0] r522;
        reg [31:0] r523;
        reg [1152:0] r524;
        reg [511:0] r525;
        reg [31:0] r526;
        reg [1152:0] r527;
        reg [511:0] r528;
        reg [31:0] r529;
        reg [1152:0] r530;
        reg [1152:0] r531;
        reg [1152:0] r532;
        reg [640:0] r533;
        reg [0:0] r534;
        reg [0:0] r536;
        reg [1153:0] r537;
        reg [1:0] r538;
        reg [27:0] r539;
        reg [41:0] r540;
        reg [34:0] r541;
        reg [20:0] r542;
        reg [48:0] r543;
        reg [50:0] r544;
        reg [38:0] r545;
        reg [49:0] r546;
        reg [37:0] r547;
        reg [42:0] r548;
        reg [56:0] r549;
        reg [33:0] r550;
        reg [44:0] r551;
        reg [53:0] r552;
        reg [16:0] r553;
        reg [18:0] r554;
        reg [6:0] r555;
        reg [17:0] r556;
        reg [5:0] r557;
        reg [10:0] r558;
        reg [24:0] r559;
        reg [1:0] r560;
        reg [12:0] r561;
        reg [21:0] r562;
        localparam l0 = 1153'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011011111000001100110100011001000111111000001111011001101010111001101100000101011010001000110001010001000011100101001001111111101001010100111111110101001110100011110001101110111100110111001010111011011001111010111010000101011010100000100111100110011001110101101111100000110011010001100100011111100000111101100110101011100110110000010101101000100011000101000100001110010100100111111110100101010011111111010100111010001111000110111011110011011100101011101101100111101011101000010101101010000010011110011001100111;
        localparam l1 = 1153'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
        localparam l2 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000;
        localparam l3 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000;
        localparam l18 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000;
        localparam l19 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000;
        localparam l20 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
        localparam l21 = 64'b0000000000000000000000000000000000000000000000000000000000000001;
        localparam l22 = 64'b0000000000000000000000000000000000000000000000000000000000000010;
        localparam l23 = 64'b0000000000000000000000000000000000000000000000000000000000000011;
        localparam l24 = 64'b0000000000000000000000000000000000000000000000000000000000000100;
        localparam l25 = 64'b0000000000000000000000000000000000000000000000000000000000000101;
        localparam l26 = 64'b0000000000000000000000000000000000000000000000000000000000000110;
        localparam l27 = 64'b0000000000000000000000000000000000000000000000000000000000000111;
        localparam l28 = 64'b0000000000000000000000000000000000000000000000000000000000001000;
        localparam l29 = 64'b0000000000000000000000000000000000000000000000000000000000001001;
        localparam l30 = 64'b0000000000000000000000000000000000000000000000000000000000001010;
        localparam l31 = 64'b0000000000000000000000000000000000000000000000000000000000001011;
        localparam l32 = 64'b0000000000000000000000000000000000000000000000000000000000001100;
        localparam l33 = 64'b0000000000000000000000000000000000000000000000000000000000001101;
        localparam l34 = 64'b0000000000000000000000000000000000000000000000000000000000001110;
        localparam l44 = 64'b0000000000000000000000000000000000000000000000000000000001000000;
        localparam l46 = 14'b00000000000000;
        localparam l47 = 8192'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110011100010111100011110010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101111101111100110100011111101110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010010001010000011011001110101100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000101111101111111111111010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100011001100011100000010000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000010011001000011110000001010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000101001010110001101101111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011101001000111110000010111011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110100000101110011011111111001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011011100111001100101001001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010011101101100010101010010010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100100011100000011001011001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110100101100001011110010110101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001110100100001110111010011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000110111011011000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001101001001100000100010110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000110101010100000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111010000001110001101011000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011010110100110010000011000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110100011001001011101000000110010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011101101100010100011010001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000010010010111000101101110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010000001101001100110010010110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010001010111111111010001010000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010011100100010110010000101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000011100001011001001001011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111011001101010000010101011101100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100101000010100111001101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100110011100000001101000100110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100110100101100011011011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101110000110110010000100111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001111011011100001010100001010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000101001001010010110011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110010100110001101010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110101011010011110010001010001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011011100000000010111111001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010111111010110010111111111000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101100000000001100100111110010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010100000110001110001100110110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010011000001111100101000101010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011101101111100110001000110110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101110010110000101010011101110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001010011101001000010010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011011110100100101100011011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000001100101000011100110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110000011001110111000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111011111011111001000111100001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110010010011011011010011100000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000001100110111111000101110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100110111101110000000110101001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000011011110101100011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110010101111100101110101110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000110001111101110000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000110001100001011011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010100000110101101100000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110000000011110101010100110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101100011100010111101101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010001111111000001010100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010110011111000100010001111100010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100101010110110000100101101100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011101001101101011101101110100101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101101011100000011111011110011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000100110111010001001001000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000010100010100010111110011000;
        localparam l48 = 32'b00000000000000000000000000000000;
        localparam l58 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001;
        localparam l59 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111;
        localparam l60 = 1'b1;
        localparam l61 = 1'b0;
        localparam l63 = 7'b0000000;
        localparam l84 = 15'b000000000000000;
        localparam l85 = 13'b0000000000000;
        localparam l86 = 25'b0000000000000000000000000;
        localparam l87 = 14'b00000000000000;
        localparam l88 = 26'b00000000000000000000000000;
        localparam l89 = 21'b000000000000000000000;
        localparam l90 = 7'b0000000;
        localparam l91 = 30'b000000000000000000000000000000;
        localparam l92 = 19'b0000000000000000000;
        localparam l93 = 10'b0000000000;
        begin
            r538 = arg_0;
            r1 = arg_1;
            r51 = arg_2;
            // let d = D::dont_care();
            //
            // if input.start {
            //    d.state = Sha256State/* fpga_test::Sha256State */ {h: [bits(H0[0]), bits(H0[1]), bits(H0[2]), bits(H0[3]), bits(H0[4]), bits(H0[5]), bits(H0[6]), bits(H0[7]), ], round: bits(0), done: false, a: bits(H0[0]), b: bits(H0[1]), c: bits(H0[2]), d: bits(H0[3]), e: bits(H0[4]), f: bits(H0[5]), g: bits(H0[6]), h_reg: bits(H0[7]),};
            //    d.w[0] = input.block[0];
            //    d.w[1] = input.block[1];
            //    d.w[2] = input.block[2];
            //    d.w[3] = input.block[3];
            //    d.w[4] = input.block[4];
            //    d.w[5] = input.block[5];
            //    d.w[6] = input.block[6];
            //    d.w[7] = input.block[7];
            //    d.w[8] = input.block[8];
            //    d.w[9] = input.block[9];
            //    d.w[10] = input.block[10];
            //    d.w[11] = input.block[11];
            //    d.w[12] = input.block[12];
            //    d.w[13] = input.block[13];
            //    d.w[14] = input.block[14];
            //    d.w[15] = input.block[15];
            // }
            //  else if !q.state.done {
            //    let round_val = q.state.round.raw();
            //    d.state = q.state;
            //    if round_val >= 16 {
            //       d.w[0] = q.w[1];
            //       d.w[1] = q.w[2];
            //       d.w[2] = q.w[3];
            //       d.w[3] = q.w[4];
            //       d.w[4] = q.w[5];
            //       d.w[5] = q.w[6];
            //       d.w[6] = q.w[7];
            //       d.w[7] = q.w[8];
            //       d.w[8] = q.w[9];
            //       d.w[9] = q.w[10];
            //       d.w[10] = q.w[11];
            //       d.w[11] = q.w[12];
            //       d.w[12] = q.w[13];
            //       d.w[13] = q.w[14];
            //       d.w[14] = q.w[15];
            //       d.w[15] = get_w(q.state.round, q.w[0], q.w[1], q.w[9], q.w[14]);
            //    }
            //     else {
            //       d.w[0] = q.w[0];
            //       d.w[1] = q.w[1];
            //       d.w[2] = q.w[2];
            //       d.w[3] = q.w[3];
            //       d.w[4] = q.w[4];
            //       d.w[5] = q.w[5];
            //       d.w[6] = q.w[6];
            //       d.w[7] = q.w[7];
            //       d.w[8] = q.w[8];
            //       d.w[9] = q.w[9];
            //       d.w[10] = q.w[10];
            //       d.w[11] = q.w[11];
            //       d.w[12] = q.w[12];
            //       d.w[13] = q.w[13];
            //       d.w[14] = q.w[14];
            //       d.w[15] = q.w[15];
            //    }
            //
            //    if round_val < 64 {
            //       let current_w = if round_val < 16 {
            //          let idx = round_val as b64;
            //          if idx == 0 {
            //             q.w[0]
            //          }
            //           else if idx == 1 {
            //             q.w[1]
            //          }
            //           else if idx == 2 {
            //             q.w[2]
            //          }
            //           else if idx == 3 {
            //             q.w[3]
            //          }
            //           else if idx == 4 {
            //             q.w[4]
            //          }
            //           else if idx == 5 {
            //             q.w[5]
            //          }
            //           else if idx == 6 {
            //             q.w[6]
            //          }
            //           else if idx == 7 {
            //             q.w[7]
            //          }
            //           else if idx == 8 {
            //             q.w[8]
            //          }
            //           else if idx == 9 {
            //             q.w[9]
            //          }
            //           else if idx == 10 {
            //             q.w[10]
            //          }
            //           else if idx == 11 {
            //             q.w[11]
            //          }
            //           else if idx == 12 {
            //             q.w[12]
            //          }
            //           else if idx == 13 {
            //             q.w[13]
            //          }
            //           else if idx == 14 {
            //             q.w[14]
            //          }
            //           else {
            //             q.w[15]
            //          }
            //
            //       }
            //        else {
            //          d.w[15]
            //       }
            //       ;
            //       let s1 = sigma1(q.state.e);
            //       let ch_result = ch(q.state.e, q.state.f, q.state.g);
            //       let temp1 = q.state.h_reg + s1 + ch_result + get_k(q.state.round) + current_w;
            //       let s0 = sigma0(q.state.a);
            //       let maj_result = maj(q.state.a, q.state.b, q.state.c);
            //       let temp2 = s0 + maj_result;
            //       d.state.h_reg = q.state.g;
            //       d.state.g = q.state.f;
            //       d.state.f = q.state.e;
            //       d.state.e = q.state.d + temp1;
            //       d.state.d = q.state.c;
            //       d.state.c = q.state.b;
            //       d.state.b = q.state.a;
            //       d.state.a = temp1 + temp2;
            //       d.state.round = bits(round_val + 1);
            //       if round_val == 63 {
            //          d.state.h[0] = q.state.h[0] + d.state.a;
            //          d.state.h[1] = q.state.h[1] + d.state.b;
            //          d.state.h[2] = q.state.h[2] + d.state.c;
            //          d.state.h[3] = q.state.h[3] + d.state.d;
            //          d.state.h[4] = q.state.h[4] + d.state.e;
            //          d.state.h[5] = q.state.h[5] + d.state.f;
            //          d.state.h[6] = q.state.h[6] + d.state.g;
            //          d.state.h[7] = q.state.h[7] + d.state.h_reg;
            //          d.state.done = true;
            //       }
            //
            //    }
            //
            // }
            //  else {
            //    d.state = q.state;
            //    d.w[0] = q.w[0];
            //    d.w[1] = q.w[1];
            //    d.w[2] = q.w[2];
            //    d.w[3] = q.w[3];
            //    d.w[4] = q.w[4];
            //    d.w[5] = q.w[5];
            //    d.w[6] = q.w[6];
            //    d.w[7] = q.w[7];
            //    d.w[8] = q.w[8];
            //    d.w[9] = q.w[9];
            //    d.w[10] = q.w[10];
            //    d.w[11] = q.w[11];
            //    d.w[12] = q.w[12];
            //    d.w[13] = q.w[13];
            //    d.w[14] = q.w[14];
            //    d.w[15] = q.w[15];
            // }
            //
            //
            r0 = r1[512];
            // d.state = Sha256State/* fpga_test::Sha256State */ {h: [bits(H0[0]), bits(H0[1]), bits(H0[2]), bits(H0[3]), bits(H0[4]), bits(H0[5]), bits(H0[6]), bits(H0[7]), ], round: bits(0), done: false, a: bits(H0[0]), b: bits(H0[1]), c: bits(H0[2]), d: bits(H0[3]), e: bits(H0[4]), f: bits(H0[5]), g: bits(H0[6]), h_reg: bits(H0[7]),};
            //
            // d.w[0] = input.block[0];
            //
            r2 = r1[511:0];
            r3 = r2[31:0];
            r4 = l0; r4[672:641] = r3;
            // d.w[1] = input.block[1];
            //
            r5 = r1[511:0];
            r6 = r5[63:32];
            r7 = r4; r7[704:673] = r6;
            // d.w[2] = input.block[2];
            //
            r8 = r1[511:0];
            r9 = r8[95:64];
            r10 = r7; r10[736:705] = r9;
            // d.w[3] = input.block[3];
            //
            r11 = r1[511:0];
            r12 = r11[127:96];
            r13 = r10; r13[768:737] = r12;
            // d.w[4] = input.block[4];
            //
            r14 = r1[511:0];
            r15 = r14[159:128];
            r16 = r13; r16[800:769] = r15;
            // d.w[5] = input.block[5];
            //
            r17 = r1[511:0];
            r18 = r17[191:160];
            r19 = r16; r19[832:801] = r18;
            // d.w[6] = input.block[6];
            //
            r20 = r1[511:0];
            r21 = r20[223:192];
            r22 = r19; r22[864:833] = r21;
            // d.w[7] = input.block[7];
            //
            r23 = r1[511:0];
            r24 = r23[255:224];
            r25 = r22; r25[896:865] = r24;
            // d.w[8] = input.block[8];
            //
            r26 = r1[511:0];
            r27 = r26[287:256];
            r28 = r25; r28[928:897] = r27;
            // d.w[9] = input.block[9];
            //
            r29 = r1[511:0];
            r30 = r29[319:288];
            r31 = r28; r31[960:929] = r30;
            // d.w[10] = input.block[10];
            //
            r32 = r1[511:0];
            r33 = r32[351:320];
            r34 = r31; r34[992:961] = r33;
            // d.w[11] = input.block[11];
            //
            r35 = r1[511:0];
            r36 = r35[383:352];
            r37 = r34; r37[1024:993] = r36;
            // d.w[12] = input.block[12];
            //
            r38 = r1[511:0];
            r39 = r38[415:384];
            r40 = r37; r40[1056:1025] = r39;
            // d.w[13] = input.block[13];
            //
            r41 = r1[511:0];
            r42 = r41[447:416];
            r43 = r40; r43[1088:1057] = r42;
            // d.w[14] = input.block[14];
            //
            r44 = r1[511:0];
            r45 = r44[479:448];
            r46 = r43; r46[1120:1089] = r45;
            // d.w[15] = input.block[15];
            //
            r47 = r1[511:0];
            r48 = r47[511:480];
            r49 = r46; r49[1152:1121] = r48;
            r50 = r51[640:0];
            r52 = r50[640];
            r53 = ~(r52);
            // let round_val = q.state.round.raw();
            //
            r54 = r51[640:0];
            r55 = r54[639:512];
            // d.state = q.state;
            //
            r56 = r51[640:0];
            r57 = l1; r57[640:0] = r56;
            // if round_val >= 16 {
            //    d.w[0] = q.w[1];
            //    d.w[1] = q.w[2];
            //    d.w[2] = q.w[3];
            //    d.w[3] = q.w[4];
            //    d.w[4] = q.w[5];
            //    d.w[5] = q.w[6];
            //    d.w[6] = q.w[7];
            //    d.w[7] = q.w[8];
            //    d.w[8] = q.w[9];
            //    d.w[9] = q.w[10];
            //    d.w[10] = q.w[11];
            //    d.w[11] = q.w[12];
            //    d.w[12] = q.w[13];
            //    d.w[13] = q.w[14];
            //    d.w[14] = q.w[15];
            //    d.w[15] = get_w(q.state.round, q.w[0], q.w[1], q.w[9], q.w[14]);
            // }
            //  else {
            //    d.w[0] = q.w[0];
            //    d.w[1] = q.w[1];
            //    d.w[2] = q.w[2];
            //    d.w[3] = q.w[3];
            //    d.w[4] = q.w[4];
            //    d.w[5] = q.w[5];
            //    d.w[6] = q.w[6];
            //    d.w[7] = q.w[7];
            //    d.w[8] = q.w[8];
            //    d.w[9] = q.w[9];
            //    d.w[10] = q.w[10];
            //    d.w[11] = q.w[11];
            //    d.w[12] = q.w[12];
            //    d.w[13] = q.w[13];
            //    d.w[14] = q.w[14];
            //    d.w[15] = q.w[15];
            // }
            //
            //
            r58 = r55 >= l2;
            // d.w[0] = q.w[1];
            //
            r59 = r51[1152:641];
            r60 = r59[63:32];
            r61 = r57; r61[672:641] = r60;
            // d.w[1] = q.w[2];
            //
            r62 = r51[1152:641];
            r63 = r62[95:64];
            r64 = r61; r64[704:673] = r63;
            // d.w[2] = q.w[3];
            //
            r65 = r51[1152:641];
            r66 = r65[127:96];
            r67 = r64; r67[736:705] = r66;
            // d.w[3] = q.w[4];
            //
            r68 = r51[1152:641];
            r69 = r68[159:128];
            r70 = r67; r70[768:737] = r69;
            // d.w[4] = q.w[5];
            //
            r71 = r51[1152:641];
            r72 = r71[191:160];
            r73 = r70; r73[800:769] = r72;
            // d.w[5] = q.w[6];
            //
            r74 = r51[1152:641];
            r75 = r74[223:192];
            r76 = r73; r76[832:801] = r75;
            // d.w[6] = q.w[7];
            //
            r77 = r51[1152:641];
            r78 = r77[255:224];
            r79 = r76; r79[864:833] = r78;
            // d.w[7] = q.w[8];
            //
            r80 = r51[1152:641];
            r81 = r80[287:256];
            r82 = r79; r82[896:865] = r81;
            // d.w[8] = q.w[9];
            //
            r83 = r51[1152:641];
            r84 = r83[319:288];
            r85 = r82; r85[928:897] = r84;
            // d.w[9] = q.w[10];
            //
            r86 = r51[1152:641];
            r87 = r86[351:320];
            r88 = r85; r88[960:929] = r87;
            // d.w[10] = q.w[11];
            //
            r89 = r51[1152:641];
            r90 = r89[383:352];
            r91 = r88; r91[992:961] = r90;
            // d.w[11] = q.w[12];
            //
            r92 = r51[1152:641];
            r93 = r92[415:384];
            r94 = r91; r94[1024:993] = r93;
            // d.w[12] = q.w[13];
            //
            r95 = r51[1152:641];
            r96 = r95[447:416];
            r97 = r94; r97[1056:1025] = r96;
            // d.w[13] = q.w[14];
            //
            r98 = r51[1152:641];
            r99 = r98[479:448];
            r100 = r97; r100[1088:1057] = r99;
            // d.w[14] = q.w[15];
            //
            r101 = r51[1152:641];
            r102 = r101[511:480];
            r103 = r100; r103[1120:1089] = r102;
            // d.w[15] = get_w(q.state.round, q.w[0], q.w[1], q.w[9], q.w[14]);
            //
            r104 = r51[640:0];
            r105 = r104[639:512];
            r106 = r51[1152:641];
            r107 = r106[31:0];
            r108 = r51[1152:641];
            r109 = r108[63:32];
            r110 = r51[1152:641];
            r111 = r110[319:288];
            r112 = r51[1152:641];
            r113 = r112[479:448];
            // let r = round.raw();
            //
            // if r < 16 {
            //    w0
            // }
            //  else {
            //    gamma1(w14) + w9 + gamma0(w1) + w0
            // }
            //
            //
            r120 = r105 < l3;
            // w0
            //
            // gamma1(w14) + w9 + gamma0(w1) + w0
            //
            // rotr(x, 17) ^ rotr(x, 19) ^ (x >> 10)
            //
            // let n = n & 31;
            //
            // (x >> n) | (x << (32 - n))
            //
            r543 = { {17{1'b0}}, r113 };
            r125 = r543[48:17];
            r553 = r113[16:0];
            r127 = { r553, l84 };
            r128 = r125 | r127;
            // let n = n & 31;
            //
            // (x >> n) | (x << (32 - n))
            //
            r544 = { {19{1'b0}}, r113 };
            r133 = r544[50:19];
            r554 = r113[18:0];
            r135 = { r554, l85 };
            r136 = r133 | r135;
            r138 = r128 ^ r136;
            r540 = { {10{1'b0}}, r113 };
            r139 = r540[41:10];
            r140 = r138 ^ r139;
            r142 = r140 + r111;
            // rotr(x, 7) ^ rotr(x, 18) ^ (x >> 3)
            //
            // let n = n & 31;
            //
            // (x >> n) | (x << (32 - n))
            //
            r545 = { {7{1'b0}}, r109 };
            r147 = r545[38:7];
            r555 = r109[6:0];
            r149 = { r555, l86 };
            r150 = r147 | r149;
            // let n = n & 31;
            //
            // (x >> n) | (x << (32 - n))
            //
            r546 = { {18{1'b0}}, r109 };
            r155 = r546[49:18];
            r556 = r109[17:0];
            r157 = { r556, l87 };
            r158 = r155 | r157;
            r160 = r150 ^ r158;
            r541 = { {3{1'b0}}, r109 };
            r161 = r541[34:3];
            r162 = r160 ^ r161;
            r164 = r142 + r162;
            r165 = r164 + r107;
            r119 = (r120) ? (r107) : (r165);
            r167 = r103; r167[1152:1121] = r119;
            // d.w[0] = q.w[0];
            //
            r168 = r51[1152:641];
            r169 = r168[31:0];
            r170 = r57; r170[672:641] = r169;
            // d.w[1] = q.w[1];
            //
            r171 = r51[1152:641];
            r172 = r171[63:32];
            r173 = r170; r173[704:673] = r172;
            // d.w[2] = q.w[2];
            //
            r174 = r51[1152:641];
            r175 = r174[95:64];
            r176 = r173; r176[736:705] = r175;
            // d.w[3] = q.w[3];
            //
            r177 = r51[1152:641];
            r178 = r177[127:96];
            r179 = r176; r179[768:737] = r178;
            // d.w[4] = q.w[4];
            //
            r180 = r51[1152:641];
            r181 = r180[159:128];
            r182 = r179; r182[800:769] = r181;
            // d.w[5] = q.w[5];
            //
            r183 = r51[1152:641];
            r184 = r183[191:160];
            r185 = r182; r185[832:801] = r184;
            // d.w[6] = q.w[6];
            //
            r186 = r51[1152:641];
            r187 = r186[223:192];
            r188 = r185; r188[864:833] = r187;
            // d.w[7] = q.w[7];
            //
            r189 = r51[1152:641];
            r190 = r189[255:224];
            r191 = r188; r191[896:865] = r190;
            // d.w[8] = q.w[8];
            //
            r192 = r51[1152:641];
            r193 = r192[287:256];
            r194 = r191; r194[928:897] = r193;
            // d.w[9] = q.w[9];
            //
            r195 = r51[1152:641];
            r196 = r195[319:288];
            r197 = r194; r197[960:929] = r196;
            // d.w[10] = q.w[10];
            //
            r198 = r51[1152:641];
            r199 = r198[351:320];
            r200 = r197; r200[992:961] = r199;
            // d.w[11] = q.w[11];
            //
            r201 = r51[1152:641];
            r202 = r201[383:352];
            r203 = r200; r203[1024:993] = r202;
            // d.w[12] = q.w[12];
            //
            r204 = r51[1152:641];
            r205 = r204[415:384];
            r206 = r203; r206[1056:1025] = r205;
            // d.w[13] = q.w[13];
            //
            r207 = r51[1152:641];
            r208 = r207[447:416];
            r209 = r206; r209[1088:1057] = r208;
            // d.w[14] = q.w[14];
            //
            r210 = r51[1152:641];
            r211 = r210[479:448];
            r212 = r209; r212[1120:1089] = r211;
            // d.w[15] = q.w[15];
            //
            r213 = r51[1152:641];
            r214 = r213[511:480];
            r215 = r212; r215[1152:1121] = r214;
            r216 = (r58) ? (r167) : (r215);
            // if round_val < 64 {
            //    let current_w = if round_val < 16 {
            //       let idx = round_val as b64;
            //       if idx == 0 {
            //          q.w[0]
            //       }
            //        else if idx == 1 {
            //          q.w[1]
            //       }
            //        else if idx == 2 {
            //          q.w[2]
            //       }
            //        else if idx == 3 {
            //          q.w[3]
            //       }
            //        else if idx == 4 {
            //          q.w[4]
            //       }
            //        else if idx == 5 {
            //          q.w[5]
            //       }
            //        else if idx == 6 {
            //          q.w[6]
            //       }
            //        else if idx == 7 {
            //          q.w[7]
            //       }
            //        else if idx == 8 {
            //          q.w[8]
            //       }
            //        else if idx == 9 {
            //          q.w[9]
            //       }
            //        else if idx == 10 {
            //          q.w[10]
            //       }
            //        else if idx == 11 {
            //          q.w[11]
            //       }
            //        else if idx == 12 {
            //          q.w[12]
            //       }
            //        else if idx == 13 {
            //          q.w[13]
            //       }
            //        else if idx == 14 {
            //          q.w[14]
            //       }
            //        else {
            //          q.w[15]
            //       }
            //
            //    }
            //     else {
            //       d.w[15]
            //    }
            //    ;
            //    let s1 = sigma1(q.state.e);
            //    let ch_result = ch(q.state.e, q.state.f, q.state.g);
            //    let temp1 = q.state.h_reg + s1 + ch_result + get_k(q.state.round) + current_w;
            //    let s0 = sigma0(q.state.a);
            //    let maj_result = maj(q.state.a, q.state.b, q.state.c);
            //    let temp2 = s0 + maj_result;
            //    d.state.h_reg = q.state.g;
            //    d.state.g = q.state.f;
            //    d.state.f = q.state.e;
            //    d.state.e = q.state.d + temp1;
            //    d.state.d = q.state.c;
            //    d.state.c = q.state.b;
            //    d.state.b = q.state.a;
            //    d.state.a = temp1 + temp2;
            //    d.state.round = bits(round_val + 1);
            //    if round_val == 63 {
            //       d.state.h[0] = q.state.h[0] + d.state.a;
            //       d.state.h[1] = q.state.h[1] + d.state.b;
            //       d.state.h[2] = q.state.h[2] + d.state.c;
            //       d.state.h[3] = q.state.h[3] + d.state.d;
            //       d.state.h[4] = q.state.h[4] + d.state.e;
            //       d.state.h[5] = q.state.h[5] + d.state.f;
            //       d.state.h[6] = q.state.h[6] + d.state.g;
            //       d.state.h[7] = q.state.h[7] + d.state.h_reg;
            //       d.state.done = true;
            //    }
            //
            // }
            //
            //
            r217 = r55 < l18;
            // let current_w = if round_val < 16 {
            //    let idx = round_val as b64;
            //    if idx == 0 {
            //       q.w[0]
            //    }
            //     else if idx == 1 {
            //       q.w[1]
            //    }
            //     else if idx == 2 {
            //       q.w[2]
            //    }
            //     else if idx == 3 {
            //       q.w[3]
            //    }
            //     else if idx == 4 {
            //       q.w[4]
            //    }
            //     else if idx == 5 {
            //       q.w[5]
            //    }
            //     else if idx == 6 {
            //       q.w[6]
            //    }
            //     else if idx == 7 {
            //       q.w[7]
            //    }
            //     else if idx == 8 {
            //       q.w[8]
            //    }
            //     else if idx == 9 {
            //       q.w[9]
            //    }
            //     else if idx == 10 {
            //       q.w[10]
            //    }
            //     else if idx == 11 {
            //       q.w[11]
            //    }
            //     else if idx == 12 {
            //       q.w[12]
            //    }
            //     else if idx == 13 {
            //       q.w[13]
            //    }
            //     else if idx == 14 {
            //       q.w[14]
            //    }
            //     else {
            //       q.w[15]
            //    }
            //
            // }
            //  else {
            //    d.w[15]
            // }
            // ;
            //
            r218 = r55 < l19;
            // let idx = round_val as b64;
            //
            r219 = r55[63:0];
            // if idx == 0 {
            //    q.w[0]
            // }
            //  else if idx == 1 {
            //    q.w[1]
            // }
            //  else if idx == 2 {
            //    q.w[2]
            // }
            //  else if idx == 3 {
            //    q.w[3]
            // }
            //  else if idx == 4 {
            //    q.w[4]
            // }
            //  else if idx == 5 {
            //    q.w[5]
            // }
            //  else if idx == 6 {
            //    q.w[6]
            // }
            //  else if idx == 7 {
            //    q.w[7]
            // }
            //  else if idx == 8 {
            //    q.w[8]
            // }
            //  else if idx == 9 {
            //    q.w[9]
            // }
            //  else if idx == 10 {
            //    q.w[10]
            // }
            //  else if idx == 11 {
            //    q.w[11]
            // }
            //  else if idx == 12 {
            //    q.w[12]
            // }
            //  else if idx == 13 {
            //    q.w[13]
            // }
            //  else if idx == 14 {
            //    q.w[14]
            // }
            //  else {
            //    q.w[15]
            // }
            //
            //
            r220 = r219 == l20;
            // q.w[0]
            //
            r221 = r51[1152:641];
            r222 = r221[31:0];
            r223 = r219 == l21;
            // q.w[1]
            //
            r224 = r51[1152:641];
            r225 = r224[63:32];
            r226 = r219 == l22;
            // q.w[2]
            //
            r227 = r51[1152:641];
            r228 = r227[95:64];
            r229 = r219 == l23;
            // q.w[3]
            //
            r230 = r51[1152:641];
            r231 = r230[127:96];
            r232 = r219 == l24;
            // q.w[4]
            //
            r233 = r51[1152:641];
            r234 = r233[159:128];
            r235 = r219 == l25;
            // q.w[5]
            //
            r236 = r51[1152:641];
            r237 = r236[191:160];
            r238 = r219 == l26;
            // q.w[6]
            //
            r239 = r51[1152:641];
            r240 = r239[223:192];
            r241 = r219 == l27;
            // q.w[7]
            //
            r242 = r51[1152:641];
            r243 = r242[255:224];
            r244 = r219 == l28;
            // q.w[8]
            //
            r245 = r51[1152:641];
            r246 = r245[287:256];
            r247 = r219 == l29;
            // q.w[9]
            //
            r248 = r51[1152:641];
            r249 = r248[319:288];
            r250 = r219 == l30;
            // q.w[10]
            //
            r251 = r51[1152:641];
            r252 = r251[351:320];
            r253 = r219 == l31;
            // q.w[11]
            //
            r254 = r51[1152:641];
            r255 = r254[383:352];
            r256 = r219 == l32;
            // q.w[12]
            //
            r257 = r51[1152:641];
            r258 = r257[415:384];
            r259 = r219 == l33;
            // q.w[13]
            //
            r260 = r51[1152:641];
            r261 = r260[447:416];
            r262 = r219 == l34;
            // q.w[14]
            //
            r263 = r51[1152:641];
            r264 = r263[479:448];
            // q.w[15]
            //
            r265 = r51[1152:641];
            r266 = r265[511:480];
            r267 = (r262) ? (r264) : (r266);
            r268 = (r259) ? (r261) : (r267);
            r269 = (r256) ? (r258) : (r268);
            r270 = (r253) ? (r255) : (r269);
            r271 = (r250) ? (r252) : (r270);
            r272 = (r247) ? (r249) : (r271);
            r273 = (r244) ? (r246) : (r272);
            r274 = (r241) ? (r243) : (r273);
            r275 = (r238) ? (r240) : (r274);
            r276 = (r235) ? (r237) : (r275);
            r277 = (r232) ? (r234) : (r276);
            r278 = (r229) ? (r231) : (r277);
            r279 = (r226) ? (r228) : (r278);
            r280 = (r223) ? (r225) : (r279);
            r281 = (r220) ? (r222) : (r280);
            // d.w[15]
            //
            r282 = r216[1152:641];
            r283 = r282[511:480];
            r284 = (r218) ? (r281) : (r283);
            // let s1 = sigma1(q.state.e);
            //
            r285 = r51[640:0];
            r286 = r285[415:384];
            // rotr(x, 6) ^ rotr(x, 11) ^ rotr(x, 25)
            //
            // let n = n & 31;
            //
            // (x >> n) | (x << (32 - n))
            //
            r547 = { {6{1'b0}}, r286 };
            r292 = r547[37:6];
            r557 = r286[5:0];
            r294 = { r557, l88 };
            r295 = r292 | r294;
            // let n = n & 31;
            //
            // (x >> n) | (x << (32 - n))
            //
            r548 = { {11{1'b0}}, r286 };
            r300 = r548[42:11];
            r558 = r286[10:0];
            r302 = { r558, l89 };
            r303 = r300 | r302;
            r305 = r295 ^ r303;
            // let n = n & 31;
            //
            // (x >> n) | (x << (32 - n))
            //
            r549 = { {25{1'b0}}, r286 };
            r309 = r549[56:25];
            r559 = r286[24:0];
            r311 = { r559, l90 };
            r312 = r309 | r311;
            r288 = r305 ^ r312;
            // let ch_result = ch(q.state.e, q.state.f, q.state.g);
            //
            r315 = r51[640:0];
            r316 = r315[415:384];
            r317 = r51[640:0];
            r318 = r317[447:416];
            r319 = r51[640:0];
            r320 = r319[479:448];
            // (x & y) ^ (!x & z)
            //
            r325 = r316 & r318;
            r326 = ~(r316);
            r327 = r326 & r320;
            r324 = r325 ^ r327;
            // let temp1 = q.state.h_reg + s1 + ch_result + get_k(q.state.round) + current_w;
            //
            r329 = r51[640:0];
            r330 = r329[511:480];
            r331 = r330 + r288;
            r332 = r331 + r324;
            r333 = r51[640:0];
            r334 = r333[639:512];
            // let r = round.raw() as b64;
            //
            r337 = r334[63:0];
            // if r < 64 {
            //    bits(K[r])
            // }
            //  else {
            //    bits(0)
            // }
            //
            //
            r338 = r337 < l44;
            // bits(K[r])
            //
            r339 = r337[13:0];
            r539 = { {14{1'b0}}, r339 };
            r542 = r539[20:0];
            r340 = { r542, l63 };
            r341 = r340[13:0];
            r342 = l46 + r341;
            r343 = l47[(r342) +: 128];
            r344 = r343[31:0];
            // bits(0)
            //
            r336 = (r338) ? (r344) : (l48);
            r346 = r332 + r336;
            r347 = r346 + r284;
            // let s0 = sigma0(q.state.a);
            //
            r348 = r51[640:0];
            r349 = r348[287:256];
            // rotr(x, 2) ^ rotr(x, 13) ^ rotr(x, 22)
            //
            // let n = n & 31;
            //
            // (x >> n) | (x << (32 - n))
            //
            r550 = { {2{1'b0}}, r349 };
            r355 = r550[33:2];
            r560 = r349[1:0];
            r357 = { r560, l91 };
            r358 = r355 | r357;
            // let n = n & 31;
            //
            // (x >> n) | (x << (32 - n))
            //
            r551 = { {13{1'b0}}, r349 };
            r363 = r551[44:13];
            r561 = r349[12:0];
            r365 = { r561, l92 };
            r366 = r363 | r365;
            r368 = r358 ^ r366;
            // let n = n & 31;
            //
            // (x >> n) | (x << (32 - n))
            //
            r552 = { {22{1'b0}}, r349 };
            r372 = r552[53:22];
            r562 = r349[21:0];
            r374 = { r562, l93 };
            r375 = r372 | r374;
            r351 = r368 ^ r375;
            // let maj_result = maj(q.state.a, q.state.b, q.state.c);
            //
            r378 = r51[640:0];
            r379 = r378[287:256];
            r380 = r51[640:0];
            r381 = r380[319:288];
            r382 = r51[640:0];
            r383 = r382[351:320];
            // (x & y) ^ (x & z) ^ (y & z)
            //
            r388 = r379 & r381;
            r389 = r379 & r383;
            r390 = r388 ^ r389;
            r391 = r381 & r383;
            r387 = r390 ^ r391;
            // let temp2 = s0 + maj_result;
            //
            r393 = r351 + r387;
            // d.state.h_reg = q.state.g;
            //
            r394 = r51[640:0];
            r395 = r394[479:448];
            r396 = r216; r396[511:480] = r395;
            // d.state.g = q.state.f;
            //
            r397 = r51[640:0];
            r398 = r397[447:416];
            r399 = r396; r399[479:448] = r398;
            // d.state.f = q.state.e;
            //
            r400 = r51[640:0];
            r401 = r400[415:384];
            r402 = r399; r402[447:416] = r401;
            // d.state.e = q.state.d + temp1;
            //
            r403 = r51[640:0];
            r404 = r403[383:352];
            r405 = r404 + r347;
            r406 = r402; r406[415:384] = r405;
            // d.state.d = q.state.c;
            //
            r407 = r51[640:0];
            r408 = r407[351:320];
            r409 = r406; r409[383:352] = r408;
            // d.state.c = q.state.b;
            //
            r410 = r51[640:0];
            r411 = r410[319:288];
            r412 = r409; r412[351:320] = r411;
            // d.state.b = q.state.a;
            //
            r413 = r51[640:0];
            r414 = r413[287:256];
            r415 = r412; r415[319:288] = r414;
            // d.state.a = temp1 + temp2;
            //
            r416 = r347 + r393;
            r417 = r415; r417[287:256] = r416;
            // d.state.round = bits(round_val + 1);
            //
            r418 = r55 + l58;
            r419 = r418[127:0];
            r420 = r417; r420[639:512] = r419;
            // if round_val == 63 {
            //    d.state.h[0] = q.state.h[0] + d.state.a;
            //    d.state.h[1] = q.state.h[1] + d.state.b;
            //    d.state.h[2] = q.state.h[2] + d.state.c;
            //    d.state.h[3] = q.state.h[3] + d.state.d;
            //    d.state.h[4] = q.state.h[4] + d.state.e;
            //    d.state.h[5] = q.state.h[5] + d.state.f;
            //    d.state.h[6] = q.state.h[6] + d.state.g;
            //    d.state.h[7] = q.state.h[7] + d.state.h_reg;
            //    d.state.done = true;
            // }
            //
            //
            r421 = r55 == l59;
            // d.state.h[0] = q.state.h[0] + d.state.a;
            //
            r422 = r51[640:0];
            r423 = r422[255:0];
            r424 = r423[31:0];
            r425 = r420[640:0];
            r426 = r425[287:256];
            r427 = r424 + r426;
            r428 = r420; r428[31:0] = r427;
            // d.state.h[1] = q.state.h[1] + d.state.b;
            //
            r429 = r51[640:0];
            r430 = r429[255:0];
            r431 = r430[63:32];
            r432 = r428[640:0];
            r433 = r432[319:288];
            r434 = r431 + r433;
            r435 = r428; r435[63:32] = r434;
            // d.state.h[2] = q.state.h[2] + d.state.c;
            //
            r436 = r51[640:0];
            r437 = r436[255:0];
            r438 = r437[95:64];
            r439 = r435[640:0];
            r440 = r439[351:320];
            r441 = r438 + r440;
            r442 = r435; r442[95:64] = r441;
            // d.state.h[3] = q.state.h[3] + d.state.d;
            //
            r443 = r51[640:0];
            r444 = r443[255:0];
            r445 = r444[127:96];
            r446 = r442[640:0];
            r447 = r446[383:352];
            r448 = r445 + r447;
            r449 = r442; r449[127:96] = r448;
            // d.state.h[4] = q.state.h[4] + d.state.e;
            //
            r450 = r51[640:0];
            r451 = r450[255:0];
            r452 = r451[159:128];
            r453 = r449[640:0];
            r454 = r453[415:384];
            r455 = r452 + r454;
            r456 = r449; r456[159:128] = r455;
            // d.state.h[5] = q.state.h[5] + d.state.f;
            //
            r457 = r51[640:0];
            r458 = r457[255:0];
            r459 = r458[191:160];
            r460 = r456[640:0];
            r461 = r460[447:416];
            r462 = r459 + r461;
            r463 = r456; r463[191:160] = r462;
            // d.state.h[6] = q.state.h[6] + d.state.g;
            //
            r464 = r51[640:0];
            r465 = r464[255:0];
            r466 = r465[223:192];
            r467 = r463[640:0];
            r468 = r467[479:448];
            r469 = r466 + r468;
            r470 = r463; r470[223:192] = r469;
            // d.state.h[7] = q.state.h[7] + d.state.h_reg;
            //
            r471 = r51[640:0];
            r472 = r471[255:0];
            r473 = r472[255:224];
            r474 = r470[640:0];
            r475 = r474[511:480];
            r476 = r473 + r475;
            r477 = r470; r477[255:224] = r476;
            // d.state.done = true;
            //
            r478 = r477; r478[640:640] = l60;
            r479 = (r421) ? (r478) : (r420);
            r480 = (r217) ? (r479) : (r216);
            // d.state = q.state;
            //
            r481 = r51[640:0];
            r482 = l1; r482[640:0] = r481;
            // d.w[0] = q.w[0];
            //
            r483 = r51[1152:641];
            r484 = r483[31:0];
            r485 = r482; r485[672:641] = r484;
            // d.w[1] = q.w[1];
            //
            r486 = r51[1152:641];
            r487 = r486[63:32];
            r488 = r485; r488[704:673] = r487;
            // d.w[2] = q.w[2];
            //
            r489 = r51[1152:641];
            r490 = r489[95:64];
            r491 = r488; r491[736:705] = r490;
            // d.w[3] = q.w[3];
            //
            r492 = r51[1152:641];
            r493 = r492[127:96];
            r494 = r491; r494[768:737] = r493;
            // d.w[4] = q.w[4];
            //
            r495 = r51[1152:641];
            r496 = r495[159:128];
            r497 = r494; r497[800:769] = r496;
            // d.w[5] = q.w[5];
            //
            r498 = r51[1152:641];
            r499 = r498[191:160];
            r500 = r497; r500[832:801] = r499;
            // d.w[6] = q.w[6];
            //
            r501 = r51[1152:641];
            r502 = r501[223:192];
            r503 = r500; r503[864:833] = r502;
            // d.w[7] = q.w[7];
            //
            r504 = r51[1152:641];
            r505 = r504[255:224];
            r506 = r503; r506[896:865] = r505;
            // d.w[8] = q.w[8];
            //
            r507 = r51[1152:641];
            r508 = r507[287:256];
            r509 = r506; r509[928:897] = r508;
            // d.w[9] = q.w[9];
            //
            r510 = r51[1152:641];
            r511 = r510[319:288];
            r512 = r509; r512[960:929] = r511;
            // d.w[10] = q.w[10];
            //
            r513 = r51[1152:641];
            r514 = r513[351:320];
            r515 = r512; r515[992:961] = r514;
            // d.w[11] = q.w[11];
            //
            r516 = r51[1152:641];
            r517 = r516[383:352];
            r518 = r515; r518[1024:993] = r517;
            // d.w[12] = q.w[12];
            //
            r519 = r51[1152:641];
            r520 = r519[415:384];
            r521 = r518; r521[1056:1025] = r520;
            // d.w[13] = q.w[13];
            //
            r522 = r51[1152:641];
            r523 = r522[447:416];
            r524 = r521; r524[1088:1057] = r523;
            // d.w[14] = q.w[14];
            //
            r525 = r51[1152:641];
            r526 = r525[479:448];
            r527 = r524; r527[1120:1089] = r526;
            // d.w[15] = q.w[15];
            //
            r528 = r51[1152:641];
            r529 = r528[511:480];
            r530 = r527; r530[1152:1121] = r529;
            r531 = (r53) ? (r480) : (r530);
            r532 = (r0) ? (r49) : (r531);
            // let output = Sha256Output/* fpga_test::Sha256Output */ {done: q.state.done,};
            //
            r533 = r51[640:0];
            r534 = r533[640];
            r536 = l61; r536[0:0] = r534;
            // (output, d, )
            //
            r537 = { r532, r536 };
            kernel_kernel = r537;
        end
    endfunction
endmodule
//
module top_state(input wire [1:0] clock_reset, input wire [640:0] i, output reg [640:0] o);
    wire [0:0] clock;
    wire [0:0] reset;
    initial begin
        o = 641'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    assign clock = clock_reset[0];
    assign reset = clock_reset[1];
    always @(posedge clock) begin
        if (reset)
        begin
            o <= 641'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        end else begin
            o <= i;
        end
    end
endmodule
// array of 16 x Positive edge triggered DFF holding value of type b32, with reset value of 0_b32
module top_w(input wire [1:0] clock_reset, input wire [511:0] i, output wire [511:0] o);
    top_w_0 c0 (.clock_reset(clock_reset),.i(i[31:0]),.o(o[31:0]));
    top_w_1 c1 (.clock_reset(clock_reset),.i(i[63:32]),.o(o[63:32]));
    top_w_10 c2 (.clock_reset(clock_reset),.i(i[95:64]),.o(o[95:64]));
    top_w_11 c3 (.clock_reset(clock_reset),.i(i[127:96]),.o(o[127:96]));
    top_w_12 c4 (.clock_reset(clock_reset),.i(i[159:128]),.o(o[159:128]));
    top_w_13 c5 (.clock_reset(clock_reset),.i(i[191:160]),.o(o[191:160]));
    top_w_14 c6 (.clock_reset(clock_reset),.i(i[223:192]),.o(o[223:192]));
    top_w_15 c7 (.clock_reset(clock_reset),.i(i[255:224]),.o(o[255:224]));
    top_w_2 c8 (.clock_reset(clock_reset),.i(i[287:256]),.o(o[287:256]));
    top_w_3 c9 (.clock_reset(clock_reset),.i(i[319:288]),.o(o[319:288]));
    top_w_4 c10 (.clock_reset(clock_reset),.i(i[351:320]),.o(o[351:320]));
    top_w_5 c11 (.clock_reset(clock_reset),.i(i[383:352]),.o(o[383:352]));
    top_w_6 c12 (.clock_reset(clock_reset),.i(i[415:384]),.o(o[415:384]));
    top_w_7 c13 (.clock_reset(clock_reset),.i(i[447:416]),.o(o[447:416]));
    top_w_8 c14 (.clock_reset(clock_reset),.i(i[479:448]),.o(o[479:448]));
    top_w_9 c15 (.clock_reset(clock_reset),.i(i[511:480]),.o(o[511:480]));
endmodule
//
module top_w_0(input wire [1:0] clock_reset, input wire [31:0] i, output reg [31:0] o);
    wire [0:0] clock;
    wire [0:0] reset;
    initial begin
        o = 32'b00000000000000000000000000000000;
    end
    assign clock = clock_reset[0];
    assign reset = clock_reset[1];
    always @(posedge clock) begin
        if (reset)
        begin
            o <= 32'b00000000000000000000000000000000;
        end else begin
            o <= i;
        end
    end
endmodule
//
module top_w_1(input wire [1:0] clock_reset, input wire [31:0] i, output reg [31:0] o);
    wire [0:0] clock;
    wire [0:0] reset;
    initial begin
        o = 32'b00000000000000000000000000000000;
    end
    assign clock = clock_reset[0];
    assign reset = clock_reset[1];
    always @(posedge clock) begin
        if (reset)
        begin
            o <= 32'b00000000000000000000000000000000;
        end else begin
            o <= i;
        end
    end
endmodule
//
module top_w_10(input wire [1:0] clock_reset, input wire [31:0] i, output reg [31:0] o);
    wire [0:0] clock;
    wire [0:0] reset;
    initial begin
        o = 32'b00000000000000000000000000000000;
    end
    assign clock = clock_reset[0];
    assign reset = clock_reset[1];
    always @(posedge clock) begin
        if (reset)
        begin
            o <= 32'b00000000000000000000000000000000;
        end else begin
            o <= i;
        end
    end
endmodule
//
module top_w_11(input wire [1:0] clock_reset, input wire [31:0] i, output reg [31:0] o);
    wire [0:0] clock;
    wire [0:0] reset;
    initial begin
        o = 32'b00000000000000000000000000000000;
    end
    assign clock = clock_reset[0];
    assign reset = clock_reset[1];
    always @(posedge clock) begin
        if (reset)
        begin
            o <= 32'b00000000000000000000000000000000;
        end else begin
            o <= i;
        end
    end
endmodule
//
module top_w_12(input wire [1:0] clock_reset, input wire [31:0] i, output reg [31:0] o);
    wire [0:0] clock;
    wire [0:0] reset;
    initial begin
        o = 32'b00000000000000000000000000000000;
    end
    assign clock = clock_reset[0];
    assign reset = clock_reset[1];
    always @(posedge clock) begin
        if (reset)
        begin
            o <= 32'b00000000000000000000000000000000;
        end else begin
            o <= i;
        end
    end
endmodule
//
module top_w_13(input wire [1:0] clock_reset, input wire [31:0] i, output reg [31:0] o);
    wire [0:0] clock;
    wire [0:0] reset;
    initial begin
        o = 32'b00000000000000000000000000000000;
    end
    assign clock = clock_reset[0];
    assign reset = clock_reset[1];
    always @(posedge clock) begin
        if (reset)
        begin
            o <= 32'b00000000000000000000000000000000;
        end else begin
            o <= i;
        end
    end
endmodule
//
module top_w_14(input wire [1:0] clock_reset, input wire [31:0] i, output reg [31:0] o);
    wire [0:0] clock;
    wire [0:0] reset;
    initial begin
        o = 32'b00000000000000000000000000000000;
    end
    assign clock = clock_reset[0];
    assign reset = clock_reset[1];
    always @(posedge clock) begin
        if (reset)
        begin
            o <= 32'b00000000000000000000000000000000;
        end else begin
            o <= i;
        end
    end
endmodule
//
module top_w_15(input wire [1:0] clock_reset, input wire [31:0] i, output reg [31:0] o);
    wire [0:0] clock;
    wire [0:0] reset;
    initial begin
        o = 32'b00000000000000000000000000000000;
    end
    assign clock = clock_reset[0];
    assign reset = clock_reset[1];
    always @(posedge clock) begin
        if (reset)
        begin
            o <= 32'b00000000000000000000000000000000;
        end else begin
            o <= i;
        end
    end
endmodule
//
module top_w_2(input wire [1:0] clock_reset, input wire [31:0] i, output reg [31:0] o);
    wire [0:0] clock;
    wire [0:0] reset;
    initial begin
        o = 32'b00000000000000000000000000000000;
    end
    assign clock = clock_reset[0];
    assign reset = clock_reset[1];
    always @(posedge clock) begin
        if (reset)
        begin
            o <= 32'b00000000000000000000000000000000;
        end else begin
            o <= i;
        end
    end
endmodule
//
module top_w_3(input wire [1:0] clock_reset, input wire [31:0] i, output reg [31:0] o);
    wire [0:0] clock;
    wire [0:0] reset;
    initial begin
        o = 32'b00000000000000000000000000000000;
    end
    assign clock = clock_reset[0];
    assign reset = clock_reset[1];
    always @(posedge clock) begin
        if (reset)
        begin
            o <= 32'b00000000000000000000000000000000;
        end else begin
            o <= i;
        end
    end
endmodule
//
module top_w_4(input wire [1:0] clock_reset, input wire [31:0] i, output reg [31:0] o);
    wire [0:0] clock;
    wire [0:0] reset;
    initial begin
        o = 32'b00000000000000000000000000000000;
    end
    assign clock = clock_reset[0];
    assign reset = clock_reset[1];
    always @(posedge clock) begin
        if (reset)
        begin
            o <= 32'b00000000000000000000000000000000;
        end else begin
            o <= i;
        end
    end
endmodule
//
module top_w_5(input wire [1:0] clock_reset, input wire [31:0] i, output reg [31:0] o);
    wire [0:0] clock;
    wire [0:0] reset;
    initial begin
        o = 32'b00000000000000000000000000000000;
    end
    assign clock = clock_reset[0];
    assign reset = clock_reset[1];
    always @(posedge clock) begin
        if (reset)
        begin
            o <= 32'b00000000000000000000000000000000;
        end else begin
            o <= i;
        end
    end
endmodule
//
module top_w_6(input wire [1:0] clock_reset, input wire [31:0] i, output reg [31:0] o);
    wire [0:0] clock;
    wire [0:0] reset;
    initial begin
        o = 32'b00000000000000000000000000000000;
    end
    assign clock = clock_reset[0];
    assign reset = clock_reset[1];
    always @(posedge clock) begin
        if (reset)
        begin
            o <= 32'b00000000000000000000000000000000;
        end else begin
            o <= i;
        end
    end
endmodule
//
module top_w_7(input wire [1:0] clock_reset, input wire [31:0] i, output reg [31:0] o);
    wire [0:0] clock;
    wire [0:0] reset;
    initial begin
        o = 32'b00000000000000000000000000000000;
    end
    assign clock = clock_reset[0];
    assign reset = clock_reset[1];
    always @(posedge clock) begin
        if (reset)
        begin
            o <= 32'b00000000000000000000000000000000;
        end else begin
            o <= i;
        end
    end
endmodule
//
module top_w_8(input wire [1:0] clock_reset, input wire [31:0] i, output reg [31:0] o);
    wire [0:0] clock;
    wire [0:0] reset;
    initial begin
        o = 32'b00000000000000000000000000000000;
    end
    assign clock = clock_reset[0];
    assign reset = clock_reset[1];
    always @(posedge clock) begin
        if (reset)
        begin
            o <= 32'b00000000000000000000000000000000;
        end else begin
            o <= i;
        end
    end
endmodule
//
module top_w_9(input wire [1:0] clock_reset, input wire [31:0] i, output reg [31:0] o);
    wire [0:0] clock;
    wire [0:0] reset;
    initial begin
        o = 32'b00000000000000000000000000000000;
    end
    assign clock = clock_reset[0];
    assign reset = clock_reset[1];
    always @(posedge clock) begin
        if (reset)
        begin
            o <= 32'b00000000000000000000000000000000;
        end else begin
            o <= i;
        end
    end
endmodule
