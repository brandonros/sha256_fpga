// synchronous circuit fpga_test::Sha256Core
module top(input wire [1:0] clock_reset, input wire [512:0] i, output wire [256:0] o);
    wire [1409:0] od;
    wire [1152:0] d;
    wire [1152:0] q;
    assign o = od[256:0];
    top_state c0 (.clock_reset(clock_reset),.i(d[640:0]),.o(q[640:0]));
    top_w c1 (.clock_reset(clock_reset),.i(d[1152:641]),.o(q[1152:641]));
    assign od = kernel_kernel(clock_reset, i, q);
    assign d = od[1409:257];
    function [1409:0] kernel_kernel(input reg [1:0] arg_0, input reg [512:0] arg_1, input reg [1152:0] arg_2);
        reg [640:0] r0;
        reg [1152:0] r1;
        reg [255:0] r2;
        reg [0:0] r3;
        reg [512:0] r4;
        reg [511:0] r5;
        reg [31:0] r6;
        reg [1152:0] r7;
        reg [511:0] r8;
        reg [31:0] r9;
        reg [1152:0] r10;
        reg [511:0] r11;
        reg [31:0] r12;
        reg [1152:0] r13;
        reg [511:0] r14;
        reg [31:0] r15;
        reg [1152:0] r16;
        reg [511:0] r17;
        reg [31:0] r18;
        reg [1152:0] r19;
        reg [511:0] r20;
        reg [31:0] r21;
        reg [1152:0] r22;
        reg [511:0] r23;
        reg [31:0] r24;
        reg [1152:0] r25;
        reg [511:0] r26;
        reg [31:0] r27;
        reg [1152:0] r28;
        reg [511:0] r29;
        reg [31:0] r30;
        reg [1152:0] r31;
        reg [511:0] r32;
        reg [31:0] r33;
        reg [1152:0] r34;
        reg [511:0] r35;
        reg [31:0] r36;
        reg [1152:0] r37;
        reg [511:0] r38;
        reg [31:0] r39;
        reg [1152:0] r40;
        reg [511:0] r41;
        reg [31:0] r42;
        reg [1152:0] r43;
        reg [511:0] r44;
        reg [31:0] r45;
        reg [1152:0] r46;
        reg [511:0] r47;
        reg [31:0] r48;
        reg [1152:0] r49;
        reg [511:0] r50;
        reg [31:0] r51;
        reg [1152:0] r52;
        reg [640:0] r53;
        reg [0:0] r54;
        reg [0:0] r55;
        reg [640:0] r56;
        reg [127:0] r57;
        reg [640:0] r58;
        reg [1152:0] r59;
        reg [0:0] r60;
        reg [511:0] r61;
        reg [31:0] r62;
        reg [1152:0] r63;
        reg [511:0] r64;
        reg [31:0] r65;
        reg [1152:0] r66;
        reg [511:0] r67;
        reg [31:0] r68;
        reg [1152:0] r69;
        reg [511:0] r70;
        reg [31:0] r71;
        reg [1152:0] r72;
        reg [511:0] r73;
        reg [31:0] r74;
        reg [1152:0] r75;
        reg [511:0] r76;
        reg [31:0] r77;
        reg [1152:0] r78;
        reg [511:0] r79;
        reg [31:0] r80;
        reg [1152:0] r81;
        reg [511:0] r82;
        reg [31:0] r83;
        reg [1152:0] r84;
        reg [511:0] r85;
        reg [31:0] r86;
        reg [1152:0] r87;
        reg [511:0] r88;
        reg [31:0] r89;
        reg [1152:0] r90;
        reg [511:0] r91;
        reg [31:0] r92;
        reg [1152:0] r93;
        reg [511:0] r94;
        reg [31:0] r95;
        reg [1152:0] r96;
        reg [511:0] r97;
        reg [31:0] r98;
        reg [1152:0] r99;
        reg [511:0] r100;
        reg [31:0] r101;
        reg [1152:0] r102;
        reg [511:0] r103;
        reg [31:0] r104;
        reg [1152:0] r105;
        reg [640:0] r106;
        reg [127:0] r107;
        reg [511:0] r108;
        reg [31:0] r109;
        reg [511:0] r110;
        reg [31:0] r111;
        reg [511:0] r112;
        reg [31:0] r113;
        reg [511:0] r114;
        reg [31:0] r115;
        reg [31:0] r121;
        reg [0:0] r122;
        reg [31:0] r127;
        reg [31:0] r129;
        reg [31:0] r130;
        reg [31:0] r135;
        reg [31:0] r137;
        reg [31:0] r138;
        reg [31:0] r140;
        reg [31:0] r141;
        reg [31:0] r142;
        reg [31:0] r144;
        reg [31:0] r149;
        reg [31:0] r151;
        reg [31:0] r152;
        reg [31:0] r157;
        reg [31:0] r159;
        reg [31:0] r160;
        reg [31:0] r162;
        reg [31:0] r163;
        reg [31:0] r164;
        reg [31:0] r166;
        reg [31:0] r167;
        reg [1152:0] r169;
        reg [511:0] r170;
        reg [31:0] r171;
        reg [1152:0] r172;
        reg [511:0] r173;
        reg [31:0] r174;
        reg [1152:0] r175;
        reg [511:0] r176;
        reg [31:0] r177;
        reg [1152:0] r178;
        reg [511:0] r179;
        reg [31:0] r180;
        reg [1152:0] r181;
        reg [511:0] r182;
        reg [31:0] r183;
        reg [1152:0] r184;
        reg [511:0] r185;
        reg [31:0] r186;
        reg [1152:0] r187;
        reg [511:0] r188;
        reg [31:0] r189;
        reg [1152:0] r190;
        reg [511:0] r191;
        reg [31:0] r192;
        reg [1152:0] r193;
        reg [511:0] r194;
        reg [31:0] r195;
        reg [1152:0] r196;
        reg [511:0] r197;
        reg [31:0] r198;
        reg [1152:0] r199;
        reg [511:0] r200;
        reg [31:0] r201;
        reg [1152:0] r202;
        reg [511:0] r203;
        reg [31:0] r204;
        reg [1152:0] r205;
        reg [511:0] r206;
        reg [31:0] r207;
        reg [1152:0] r208;
        reg [511:0] r209;
        reg [31:0] r210;
        reg [1152:0] r211;
        reg [511:0] r212;
        reg [31:0] r213;
        reg [1152:0] r214;
        reg [511:0] r215;
        reg [31:0] r216;
        reg [1152:0] r217;
        reg [1152:0] r218;
        reg [0:0] r219;
        reg [0:0] r220;
        reg [63:0] r221;
        reg [0:0] r222;
        reg [511:0] r223;
        reg [31:0] r224;
        reg [0:0] r225;
        reg [511:0] r226;
        reg [31:0] r227;
        reg [0:0] r228;
        reg [511:0] r229;
        reg [31:0] r230;
        reg [0:0] r231;
        reg [511:0] r232;
        reg [31:0] r233;
        reg [0:0] r234;
        reg [511:0] r235;
        reg [31:0] r236;
        reg [0:0] r237;
        reg [511:0] r238;
        reg [31:0] r239;
        reg [0:0] r240;
        reg [511:0] r241;
        reg [31:0] r242;
        reg [0:0] r243;
        reg [511:0] r244;
        reg [31:0] r245;
        reg [0:0] r246;
        reg [511:0] r247;
        reg [31:0] r248;
        reg [0:0] r249;
        reg [511:0] r250;
        reg [31:0] r251;
        reg [0:0] r252;
        reg [511:0] r253;
        reg [31:0] r254;
        reg [0:0] r255;
        reg [511:0] r256;
        reg [31:0] r257;
        reg [0:0] r258;
        reg [511:0] r259;
        reg [31:0] r260;
        reg [0:0] r261;
        reg [511:0] r262;
        reg [31:0] r263;
        reg [0:0] r264;
        reg [511:0] r265;
        reg [31:0] r266;
        reg [511:0] r267;
        reg [31:0] r268;
        reg [31:0] r269;
        reg [31:0] r270;
        reg [31:0] r271;
        reg [31:0] r272;
        reg [31:0] r273;
        reg [31:0] r274;
        reg [31:0] r275;
        reg [31:0] r276;
        reg [31:0] r277;
        reg [31:0] r278;
        reg [31:0] r279;
        reg [31:0] r280;
        reg [31:0] r281;
        reg [31:0] r282;
        reg [31:0] r283;
        reg [511:0] r284;
        reg [31:0] r285;
        reg [31:0] r286;
        reg [640:0] r287;
        reg [31:0] r288;
        reg [31:0] r290;
        reg [31:0] r294;
        reg [31:0] r296;
        reg [31:0] r297;
        reg [31:0] r302;
        reg [31:0] r304;
        reg [31:0] r305;
        reg [31:0] r307;
        reg [31:0] r311;
        reg [31:0] r313;
        reg [31:0] r314;
        reg [640:0] r317;
        reg [31:0] r318;
        reg [640:0] r319;
        reg [31:0] r320;
        reg [640:0] r321;
        reg [31:0] r322;
        reg [31:0] r326;
        reg [31:0] r327;
        reg [31:0] r328;
        reg [31:0] r329;
        reg [640:0] r331;
        reg [31:0] r332;
        reg [31:0] r333;
        reg [31:0] r334;
        reg [640:0] r335;
        reg [127:0] r336;
        reg [31:0] r338;
        reg [63:0] r339;
        reg [0:0] r340;
        reg [13:0] r341;
        reg [27:0] r342;
        reg [13:0] r343;
        reg [13:0] r344;
        reg [127:0] r345;
        reg [31:0] r346;
        reg [31:0] r348;
        reg [31:0] r349;
        reg [640:0] r350;
        reg [31:0] r351;
        reg [31:0] r353;
        reg [31:0] r357;
        reg [31:0] r359;
        reg [31:0] r360;
        reg [31:0] r365;
        reg [31:0] r367;
        reg [31:0] r368;
        reg [31:0] r370;
        reg [31:0] r374;
        reg [31:0] r376;
        reg [31:0] r377;
        reg [640:0] r380;
        reg [31:0] r381;
        reg [640:0] r382;
        reg [31:0] r383;
        reg [640:0] r384;
        reg [31:0] r385;
        reg [31:0] r389;
        reg [31:0] r390;
        reg [31:0] r391;
        reg [31:0] r392;
        reg [31:0] r393;
        reg [31:0] r395;
        reg [640:0] r396;
        reg [31:0] r397;
        reg [1152:0] r398;
        reg [640:0] r399;
        reg [31:0] r400;
        reg [1152:0] r401;
        reg [640:0] r402;
        reg [31:0] r403;
        reg [1152:0] r404;
        reg [640:0] r405;
        reg [31:0] r406;
        reg [31:0] r407;
        reg [1152:0] r408;
        reg [640:0] r409;
        reg [31:0] r410;
        reg [1152:0] r411;
        reg [640:0] r412;
        reg [31:0] r413;
        reg [1152:0] r414;
        reg [640:0] r415;
        reg [31:0] r416;
        reg [1152:0] r417;
        reg [31:0] r418;
        reg [1152:0] r419;
        reg [127:0] r420;
        reg [127:0] r421;
        reg [1152:0] r422;
        reg [0:0] r423;
        reg [640:0] r424;
        reg [255:0] r425;
        reg [31:0] r426;
        reg [640:0] r427;
        reg [31:0] r428;
        reg [31:0] r429;
        reg [1152:0] r430;
        reg [640:0] r431;
        reg [255:0] r432;
        reg [31:0] r433;
        reg [640:0] r434;
        reg [31:0] r435;
        reg [31:0] r436;
        reg [1152:0] r437;
        reg [640:0] r438;
        reg [255:0] r439;
        reg [31:0] r440;
        reg [640:0] r441;
        reg [31:0] r442;
        reg [31:0] r443;
        reg [1152:0] r444;
        reg [640:0] r445;
        reg [255:0] r446;
        reg [31:0] r447;
        reg [640:0] r448;
        reg [31:0] r449;
        reg [31:0] r450;
        reg [1152:0] r451;
        reg [640:0] r452;
        reg [255:0] r453;
        reg [31:0] r454;
        reg [640:0] r455;
        reg [31:0] r456;
        reg [31:0] r457;
        reg [1152:0] r458;
        reg [640:0] r459;
        reg [255:0] r460;
        reg [31:0] r461;
        reg [640:0] r462;
        reg [31:0] r463;
        reg [31:0] r464;
        reg [1152:0] r465;
        reg [640:0] r466;
        reg [255:0] r467;
        reg [31:0] r468;
        reg [640:0] r469;
        reg [31:0] r470;
        reg [31:0] r471;
        reg [1152:0] r472;
        reg [640:0] r473;
        reg [255:0] r474;
        reg [31:0] r475;
        reg [640:0] r476;
        reg [31:0] r477;
        reg [31:0] r478;
        reg [1152:0] r479;
        reg [1152:0] r480;
        reg [640:0] r481;
        reg [255:0] r482;
        reg [1152:0] r483;
        reg [255:0] r484;
        reg [0:0] r485;
        reg [1152:0] r486;
        reg [255:0] r487;
        reg [0:0] r488;
        reg [640:0] r489;
        reg [1152:0] r490;
        reg [511:0] r491;
        reg [31:0] r492;
        reg [1152:0] r493;
        reg [511:0] r494;
        reg [31:0] r495;
        reg [1152:0] r496;
        reg [511:0] r497;
        reg [31:0] r498;
        reg [1152:0] r499;
        reg [511:0] r500;
        reg [31:0] r501;
        reg [1152:0] r502;
        reg [511:0] r503;
        reg [31:0] r504;
        reg [1152:0] r505;
        reg [511:0] r506;
        reg [31:0] r507;
        reg [1152:0] r508;
        reg [511:0] r509;
        reg [31:0] r510;
        reg [1152:0] r511;
        reg [511:0] r512;
        reg [31:0] r513;
        reg [1152:0] r514;
        reg [511:0] r515;
        reg [31:0] r516;
        reg [1152:0] r517;
        reg [511:0] r518;
        reg [31:0] r519;
        reg [1152:0] r520;
        reg [511:0] r521;
        reg [31:0] r522;
        reg [1152:0] r523;
        reg [511:0] r524;
        reg [31:0] r525;
        reg [1152:0] r526;
        reg [511:0] r527;
        reg [31:0] r528;
        reg [1152:0] r529;
        reg [511:0] r530;
        reg [31:0] r531;
        reg [1152:0] r532;
        reg [511:0] r533;
        reg [31:0] r534;
        reg [1152:0] r535;
        reg [511:0] r536;
        reg [31:0] r537;
        reg [1152:0] r538;
        reg [640:0] r539;
        reg [255:0] r540;
        reg [1152:0] r541;
        reg [255:0] r542;
        reg [0:0] r543;
        reg [1152:0] r544;
        reg [255:0] r545;
        reg [0:0] r546;
        reg [256:0] r547;
        reg [1409:0] r548;
        reg [1:0] r549;
        reg [27:0] r550;
        reg [41:0] r551;
        reg [34:0] r552;
        reg [20:0] r553;
        reg [48:0] r554;
        reg [50:0] r555;
        reg [38:0] r556;
        reg [49:0] r557;
        reg [37:0] r558;
        reg [42:0] r559;
        reg [56:0] r560;
        reg [33:0] r561;
        reg [44:0] r562;
        reg [53:0] r563;
        reg [16:0] r564;
        reg [18:0] r565;
        reg [6:0] r566;
        reg [17:0] r567;
        reg [5:0] r568;
        reg [10:0] r569;
        reg [24:0] r570;
        reg [1:0] r571;
        reg [12:0] r572;
        reg [21:0] r573;
        localparam l0 = 1153'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011011111000001100110100011001000111111000001111011001101010111001101100000101011010001000110001010001000011100101001001111111101001010100111111110101001110100011110001101110111100110111001010111011011001111010111010000101011010100000100111100110011001110101101111100000110011010001100100011111100000111101100110101011100110110000010101101000100011000101000100001110010100100111111110100101010011111111010100111010001111000110111011110011011100101011101101100111101011101000010101101010000010011110011001100111;
        localparam l1 = 1153'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
        localparam l2 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000;
        localparam l3 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000;
        localparam l18 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000;
        localparam l19 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000;
        localparam l20 = 64'b0000000000000000000000000000000000000000000000000000000000000000;
        localparam l21 = 64'b0000000000000000000000000000000000000000000000000000000000000001;
        localparam l22 = 64'b0000000000000000000000000000000000000000000000000000000000000010;
        localparam l23 = 64'b0000000000000000000000000000000000000000000000000000000000000011;
        localparam l24 = 64'b0000000000000000000000000000000000000000000000000000000000000100;
        localparam l25 = 64'b0000000000000000000000000000000000000000000000000000000000000101;
        localparam l26 = 64'b0000000000000000000000000000000000000000000000000000000000000110;
        localparam l27 = 64'b0000000000000000000000000000000000000000000000000000000000000111;
        localparam l28 = 64'b0000000000000000000000000000000000000000000000000000000000001000;
        localparam l29 = 64'b0000000000000000000000000000000000000000000000000000000000001001;
        localparam l30 = 64'b0000000000000000000000000000000000000000000000000000000000001010;
        localparam l31 = 64'b0000000000000000000000000000000000000000000000000000000000001011;
        localparam l32 = 64'b0000000000000000000000000000000000000000000000000000000000001100;
        localparam l33 = 64'b0000000000000000000000000000000000000000000000000000000000001101;
        localparam l34 = 64'b0000000000000000000000000000000000000000000000000000000000001110;
        localparam l44 = 64'b0000000000000000000000000000000000000000000000000000000001000000;
        localparam l46 = 14'b00000000000000;
        localparam l47 = 8192'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000110011100010111100011110010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101111101111100110100011111101110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010010001010000011011001110101100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000101111101111111111111010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100011001100011100000010000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000010011001000011110000001010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000101001010110001101101111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011101001000111110000010111011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110100000101110011011111111001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011011100111001100101001001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010011101101100010101010010010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100100011100000011001011001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110100101100001011110010110101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001110100100001110111010011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111000110111011011000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001101001001100000100010110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000110101010100000011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111010000001110001101011000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011010110100110010000011000100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110100011001001011101000000110010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011101101100010100011010001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000010010010111000101101110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010000001101001100110010010110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010001010111111111010001010000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010011100100010110010000101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000011100001011001001001011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111011001101010000010101011101100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100101000010100111001101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010100110011100000001101000100110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100110100101100011011011111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101110000110110010000100111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001111011011100001010100001010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000101001001010010110011100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110010100110001101010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110101011010011110010001010001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100011011100000000010111111001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010111111010110010111111111000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101100000000001100100111110010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010100000110001110001100110110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010011000001111100101000101010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011101101111100110001000110110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101110010110000101010011101110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001010011101001000010010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001011011110100100101100011011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000001100101000011100110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110000011001110111000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111011111011111001000111100001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110010010011011011010011100000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000001100110111111000101110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100110111101110000000110101001110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000011011110101100011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110010101111100101110101110100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010000110001111101110000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000110001100001011011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010100000110101101100000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110000000011110101010100110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010101100011100010111101101010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010010001111111000001010100100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010110011111000100010001111100010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011100101010110110000100101101100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011101001101101011101101110100101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101101011100000011111011110011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000100110111010001001001000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000010100010100010111110011000;
        localparam l48 = 32'b00000000000000000000000000000000;
        localparam l58 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001;
        localparam l59 = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111;
        localparam l60 = 1'b1;
        localparam l61 = 1'b1;
        localparam l62 = 1'b0;
        localparam l63 = 1'b1;
        localparam l65 = 7'b0000000;
        localparam l86 = 15'b000000000000000;
        localparam l87 = 13'b0000000000000;
        localparam l88 = 25'b0000000000000000000000000;
        localparam l89 = 14'b00000000000000;
        localparam l90 = 26'b00000000000000000000000000;
        localparam l91 = 21'b000000000000000000000;
        localparam l92 = 7'b0000000;
        localparam l93 = 30'b000000000000000000000000000000;
        localparam l94 = 19'b0000000000000000000;
        localparam l95 = 10'b0000000000;
        begin
            r549 = arg_0;
            r4 = arg_1;
            r1 = arg_2;
            // let d = D::dont_care();
            //
            // let output_valid = false;
            //
            // let hash_out = q.state.h;
            //
            r0 = r1[640:0];
            r2 = r0[255:0];
            // if input.start {
            //    d.state = Sha256State/* fpga_test::Sha256State */ {h: [bits(H0[0]), bits(H0[1]), bits(H0[2]), bits(H0[3]), bits(H0[4]), bits(H0[5]), bits(H0[6]), bits(H0[7]), ], round: bits(0), done: false, a: bits(H0[0]), b: bits(H0[1]), c: bits(H0[2]), d: bits(H0[3]), e: bits(H0[4]), f: bits(H0[5]), g: bits(H0[6]), h_reg: bits(H0[7]),};
            //    d.w[0] = input.block[0];
            //    d.w[1] = input.block[1];
            //    d.w[2] = input.block[2];
            //    d.w[3] = input.block[3];
            //    d.w[4] = input.block[4];
            //    d.w[5] = input.block[5];
            //    d.w[6] = input.block[6];
            //    d.w[7] = input.block[7];
            //    d.w[8] = input.block[8];
            //    d.w[9] = input.block[9];
            //    d.w[10] = input.block[10];
            //    d.w[11] = input.block[11];
            //    d.w[12] = input.block[12];
            //    d.w[13] = input.block[13];
            //    d.w[14] = input.block[14];
            //    d.w[15] = input.block[15];
            // }
            //  else if !q.state.done {
            //    let round_val = q.state.round.raw();
            //    d.state = q.state;
            //    if round_val >= 16 {
            //       d.w[0] = q.w[1];
            //       d.w[1] = q.w[2];
            //       d.w[2] = q.w[3];
            //       d.w[3] = q.w[4];
            //       d.w[4] = q.w[5];
            //       d.w[5] = q.w[6];
            //       d.w[6] = q.w[7];
            //       d.w[7] = q.w[8];
            //       d.w[8] = q.w[9];
            //       d.w[9] = q.w[10];
            //       d.w[10] = q.w[11];
            //       d.w[11] = q.w[12];
            //       d.w[12] = q.w[13];
            //       d.w[13] = q.w[14];
            //       d.w[14] = q.w[15];
            //       d.w[15] = get_w(q.state.round, q.w[0], q.w[1], q.w[9], q.w[14]);
            //    }
            //     else {
            //       d.w[0] = q.w[0];
            //       d.w[1] = q.w[1];
            //       d.w[2] = q.w[2];
            //       d.w[3] = q.w[3];
            //       d.w[4] = q.w[4];
            //       d.w[5] = q.w[5];
            //       d.w[6] = q.w[6];
            //       d.w[7] = q.w[7];
            //       d.w[8] = q.w[8];
            //       d.w[9] = q.w[9];
            //       d.w[10] = q.w[10];
            //       d.w[11] = q.w[11];
            //       d.w[12] = q.w[12];
            //       d.w[13] = q.w[13];
            //       d.w[14] = q.w[14];
            //       d.w[15] = q.w[15];
            //    }
            //
            //    if round_val < 64 {
            //       let current_w = if round_val < 16 {
            //          let idx = round_val as b64;
            //          if idx == 0 {
            //             q.w[0]
            //          }
            //           else if idx == 1 {
            //             q.w[1]
            //          }
            //           else if idx == 2 {
            //             q.w[2]
            //          }
            //           else if idx == 3 {
            //             q.w[3]
            //          }
            //           else if idx == 4 {
            //             q.w[4]
            //          }
            //           else if idx == 5 {
            //             q.w[5]
            //          }
            //           else if idx == 6 {
            //             q.w[6]
            //          }
            //           else if idx == 7 {
            //             q.w[7]
            //          }
            //           else if idx == 8 {
            //             q.w[8]
            //          }
            //           else if idx == 9 {
            //             q.w[9]
            //          }
            //           else if idx == 10 {
            //             q.w[10]
            //          }
            //           else if idx == 11 {
            //             q.w[11]
            //          }
            //           else if idx == 12 {
            //             q.w[12]
            //          }
            //           else if idx == 13 {
            //             q.w[13]
            //          }
            //           else if idx == 14 {
            //             q.w[14]
            //          }
            //           else {
            //             q.w[15]
            //          }
            //
            //       }
            //        else {
            //          d.w[15]
            //       }
            //       ;
            //       let s1 = sigma1(q.state.e);
            //       let ch_result = ch(q.state.e, q.state.f, q.state.g);
            //       let temp1 = q.state.h_reg + s1 + ch_result + get_k(q.state.round) + current_w;
            //       let s0 = sigma0(q.state.a);
            //       let maj_result = maj(q.state.a, q.state.b, q.state.c);
            //       let temp2 = s0 + maj_result;
            //       d.state.h_reg = q.state.g;
            //       d.state.g = q.state.f;
            //       d.state.f = q.state.e;
            //       d.state.e = q.state.d + temp1;
            //       d.state.d = q.state.c;
            //       d.state.c = q.state.b;
            //       d.state.b = q.state.a;
            //       d.state.a = temp1 + temp2;
            //       d.state.round = bits(round_val + 1);
            //       if round_val == 63 {
            //          d.state.h[0] = q.state.h[0] + d.state.a;
            //          d.state.h[1] = q.state.h[1] + d.state.b;
            //          d.state.h[2] = q.state.h[2] + d.state.c;
            //          d.state.h[3] = q.state.h[3] + d.state.d;
            //          d.state.h[4] = q.state.h[4] + d.state.e;
            //          d.state.h[5] = q.state.h[5] + d.state.f;
            //          d.state.h[6] = q.state.h[6] + d.state.g;
            //          d.state.h[7] = q.state.h[7] + d.state.h_reg;
            //          d.state.done = true;
            //          output_valid = true;
            //          hash_out = d.state.h;
            //       }
            //
            //    }
            //
            // }
            //  else {
            //    d.state = q.state;
            //    d.w[0] = q.w[0];
            //    d.w[1] = q.w[1];
            //    d.w[2] = q.w[2];
            //    d.w[3] = q.w[3];
            //    d.w[4] = q.w[4];
            //    d.w[5] = q.w[5];
            //    d.w[6] = q.w[6];
            //    d.w[7] = q.w[7];
            //    d.w[8] = q.w[8];
            //    d.w[9] = q.w[9];
            //    d.w[10] = q.w[10];
            //    d.w[11] = q.w[11];
            //    d.w[12] = q.w[12];
            //    d.w[13] = q.w[13];
            //    d.w[14] = q.w[14];
            //    d.w[15] = q.w[15];
            //    output_valid = true;
            //    hash_out = q.state.h;
            // }
            //
            //
            r3 = r4[512];
            // d.state = Sha256State/* fpga_test::Sha256State */ {h: [bits(H0[0]), bits(H0[1]), bits(H0[2]), bits(H0[3]), bits(H0[4]), bits(H0[5]), bits(H0[6]), bits(H0[7]), ], round: bits(0), done: false, a: bits(H0[0]), b: bits(H0[1]), c: bits(H0[2]), d: bits(H0[3]), e: bits(H0[4]), f: bits(H0[5]), g: bits(H0[6]), h_reg: bits(H0[7]),};
            //
            // d.w[0] = input.block[0];
            //
            r5 = r4[511:0];
            r6 = r5[31:0];
            r7 = l0; r7[672:641] = r6;
            // d.w[1] = input.block[1];
            //
            r8 = r4[511:0];
            r9 = r8[63:32];
            r10 = r7; r10[704:673] = r9;
            // d.w[2] = input.block[2];
            //
            r11 = r4[511:0];
            r12 = r11[95:64];
            r13 = r10; r13[736:705] = r12;
            // d.w[3] = input.block[3];
            //
            r14 = r4[511:0];
            r15 = r14[127:96];
            r16 = r13; r16[768:737] = r15;
            // d.w[4] = input.block[4];
            //
            r17 = r4[511:0];
            r18 = r17[159:128];
            r19 = r16; r19[800:769] = r18;
            // d.w[5] = input.block[5];
            //
            r20 = r4[511:0];
            r21 = r20[191:160];
            r22 = r19; r22[832:801] = r21;
            // d.w[6] = input.block[6];
            //
            r23 = r4[511:0];
            r24 = r23[223:192];
            r25 = r22; r25[864:833] = r24;
            // d.w[7] = input.block[7];
            //
            r26 = r4[511:0];
            r27 = r26[255:224];
            r28 = r25; r28[896:865] = r27;
            // d.w[8] = input.block[8];
            //
            r29 = r4[511:0];
            r30 = r29[287:256];
            r31 = r28; r31[928:897] = r30;
            // d.w[9] = input.block[9];
            //
            r32 = r4[511:0];
            r33 = r32[319:288];
            r34 = r31; r34[960:929] = r33;
            // d.w[10] = input.block[10];
            //
            r35 = r4[511:0];
            r36 = r35[351:320];
            r37 = r34; r37[992:961] = r36;
            // d.w[11] = input.block[11];
            //
            r38 = r4[511:0];
            r39 = r38[383:352];
            r40 = r37; r40[1024:993] = r39;
            // d.w[12] = input.block[12];
            //
            r41 = r4[511:0];
            r42 = r41[415:384];
            r43 = r40; r43[1056:1025] = r42;
            // d.w[13] = input.block[13];
            //
            r44 = r4[511:0];
            r45 = r44[447:416];
            r46 = r43; r46[1088:1057] = r45;
            // d.w[14] = input.block[14];
            //
            r47 = r4[511:0];
            r48 = r47[479:448];
            r49 = r46; r49[1120:1089] = r48;
            // d.w[15] = input.block[15];
            //
            r50 = r4[511:0];
            r51 = r50[511:480];
            r52 = r49; r52[1152:1121] = r51;
            r53 = r1[640:0];
            r54 = r53[640];
            r55 = ~(r54);
            // let round_val = q.state.round.raw();
            //
            r56 = r1[640:0];
            r57 = r56[639:512];
            // d.state = q.state;
            //
            r58 = r1[640:0];
            r59 = l1; r59[640:0] = r58;
            // if round_val >= 16 {
            //    d.w[0] = q.w[1];
            //    d.w[1] = q.w[2];
            //    d.w[2] = q.w[3];
            //    d.w[3] = q.w[4];
            //    d.w[4] = q.w[5];
            //    d.w[5] = q.w[6];
            //    d.w[6] = q.w[7];
            //    d.w[7] = q.w[8];
            //    d.w[8] = q.w[9];
            //    d.w[9] = q.w[10];
            //    d.w[10] = q.w[11];
            //    d.w[11] = q.w[12];
            //    d.w[12] = q.w[13];
            //    d.w[13] = q.w[14];
            //    d.w[14] = q.w[15];
            //    d.w[15] = get_w(q.state.round, q.w[0], q.w[1], q.w[9], q.w[14]);
            // }
            //  else {
            //    d.w[0] = q.w[0];
            //    d.w[1] = q.w[1];
            //    d.w[2] = q.w[2];
            //    d.w[3] = q.w[3];
            //    d.w[4] = q.w[4];
            //    d.w[5] = q.w[5];
            //    d.w[6] = q.w[6];
            //    d.w[7] = q.w[7];
            //    d.w[8] = q.w[8];
            //    d.w[9] = q.w[9];
            //    d.w[10] = q.w[10];
            //    d.w[11] = q.w[11];
            //    d.w[12] = q.w[12];
            //    d.w[13] = q.w[13];
            //    d.w[14] = q.w[14];
            //    d.w[15] = q.w[15];
            // }
            //
            //
            r60 = r57 >= l2;
            // d.w[0] = q.w[1];
            //
            r61 = r1[1152:641];
            r62 = r61[63:32];
            r63 = r59; r63[672:641] = r62;
            // d.w[1] = q.w[2];
            //
            r64 = r1[1152:641];
            r65 = r64[95:64];
            r66 = r63; r66[704:673] = r65;
            // d.w[2] = q.w[3];
            //
            r67 = r1[1152:641];
            r68 = r67[127:96];
            r69 = r66; r69[736:705] = r68;
            // d.w[3] = q.w[4];
            //
            r70 = r1[1152:641];
            r71 = r70[159:128];
            r72 = r69; r72[768:737] = r71;
            // d.w[4] = q.w[5];
            //
            r73 = r1[1152:641];
            r74 = r73[191:160];
            r75 = r72; r75[800:769] = r74;
            // d.w[5] = q.w[6];
            //
            r76 = r1[1152:641];
            r77 = r76[223:192];
            r78 = r75; r78[832:801] = r77;
            // d.w[6] = q.w[7];
            //
            r79 = r1[1152:641];
            r80 = r79[255:224];
            r81 = r78; r81[864:833] = r80;
            // d.w[7] = q.w[8];
            //
            r82 = r1[1152:641];
            r83 = r82[287:256];
            r84 = r81; r84[896:865] = r83;
            // d.w[8] = q.w[9];
            //
            r85 = r1[1152:641];
            r86 = r85[319:288];
            r87 = r84; r87[928:897] = r86;
            // d.w[9] = q.w[10];
            //
            r88 = r1[1152:641];
            r89 = r88[351:320];
            r90 = r87; r90[960:929] = r89;
            // d.w[10] = q.w[11];
            //
            r91 = r1[1152:641];
            r92 = r91[383:352];
            r93 = r90; r93[992:961] = r92;
            // d.w[11] = q.w[12];
            //
            r94 = r1[1152:641];
            r95 = r94[415:384];
            r96 = r93; r96[1024:993] = r95;
            // d.w[12] = q.w[13];
            //
            r97 = r1[1152:641];
            r98 = r97[447:416];
            r99 = r96; r99[1056:1025] = r98;
            // d.w[13] = q.w[14];
            //
            r100 = r1[1152:641];
            r101 = r100[479:448];
            r102 = r99; r102[1088:1057] = r101;
            // d.w[14] = q.w[15];
            //
            r103 = r1[1152:641];
            r104 = r103[511:480];
            r105 = r102; r105[1120:1089] = r104;
            // d.w[15] = get_w(q.state.round, q.w[0], q.w[1], q.w[9], q.w[14]);
            //
            r106 = r1[640:0];
            r107 = r106[639:512];
            r108 = r1[1152:641];
            r109 = r108[31:0];
            r110 = r1[1152:641];
            r111 = r110[63:32];
            r112 = r1[1152:641];
            r113 = r112[319:288];
            r114 = r1[1152:641];
            r115 = r114[479:448];
            // let r = round.raw();
            //
            // if r < 16 {
            //    w0
            // }
            //  else {
            //    gamma1(w14) + w9 + gamma0(w1) + w0
            // }
            //
            //
            r122 = r107 < l3;
            // w0
            //
            // gamma1(w14) + w9 + gamma0(w1) + w0
            //
            // rotr(x, 17) ^ rotr(x, 19) ^ (x >> 10)
            //
            // let n = n & 31;
            //
            // (x >> n) | (x << (32 - n))
            //
            r554 = { {17{1'b0}}, r115 };
            r127 = r554[48:17];
            r564 = r115[16:0];
            r129 = { r564, l86 };
            r130 = r127 | r129;
            // let n = n & 31;
            //
            // (x >> n) | (x << (32 - n))
            //
            r555 = { {19{1'b0}}, r115 };
            r135 = r555[50:19];
            r565 = r115[18:0];
            r137 = { r565, l87 };
            r138 = r135 | r137;
            r140 = r130 ^ r138;
            r551 = { {10{1'b0}}, r115 };
            r141 = r551[41:10];
            r142 = r140 ^ r141;
            r144 = r142 + r113;
            // rotr(x, 7) ^ rotr(x, 18) ^ (x >> 3)
            //
            // let n = n & 31;
            //
            // (x >> n) | (x << (32 - n))
            //
            r556 = { {7{1'b0}}, r111 };
            r149 = r556[38:7];
            r566 = r111[6:0];
            r151 = { r566, l88 };
            r152 = r149 | r151;
            // let n = n & 31;
            //
            // (x >> n) | (x << (32 - n))
            //
            r557 = { {18{1'b0}}, r111 };
            r157 = r557[49:18];
            r567 = r111[17:0];
            r159 = { r567, l89 };
            r160 = r157 | r159;
            r162 = r152 ^ r160;
            r552 = { {3{1'b0}}, r111 };
            r163 = r552[34:3];
            r164 = r162 ^ r163;
            r166 = r144 + r164;
            r167 = r166 + r109;
            r121 = (r122) ? (r109) : (r167);
            r169 = r105; r169[1152:1121] = r121;
            // d.w[0] = q.w[0];
            //
            r170 = r1[1152:641];
            r171 = r170[31:0];
            r172 = r59; r172[672:641] = r171;
            // d.w[1] = q.w[1];
            //
            r173 = r1[1152:641];
            r174 = r173[63:32];
            r175 = r172; r175[704:673] = r174;
            // d.w[2] = q.w[2];
            //
            r176 = r1[1152:641];
            r177 = r176[95:64];
            r178 = r175; r178[736:705] = r177;
            // d.w[3] = q.w[3];
            //
            r179 = r1[1152:641];
            r180 = r179[127:96];
            r181 = r178; r181[768:737] = r180;
            // d.w[4] = q.w[4];
            //
            r182 = r1[1152:641];
            r183 = r182[159:128];
            r184 = r181; r184[800:769] = r183;
            // d.w[5] = q.w[5];
            //
            r185 = r1[1152:641];
            r186 = r185[191:160];
            r187 = r184; r187[832:801] = r186;
            // d.w[6] = q.w[6];
            //
            r188 = r1[1152:641];
            r189 = r188[223:192];
            r190 = r187; r190[864:833] = r189;
            // d.w[7] = q.w[7];
            //
            r191 = r1[1152:641];
            r192 = r191[255:224];
            r193 = r190; r193[896:865] = r192;
            // d.w[8] = q.w[8];
            //
            r194 = r1[1152:641];
            r195 = r194[287:256];
            r196 = r193; r196[928:897] = r195;
            // d.w[9] = q.w[9];
            //
            r197 = r1[1152:641];
            r198 = r197[319:288];
            r199 = r196; r199[960:929] = r198;
            // d.w[10] = q.w[10];
            //
            r200 = r1[1152:641];
            r201 = r200[351:320];
            r202 = r199; r202[992:961] = r201;
            // d.w[11] = q.w[11];
            //
            r203 = r1[1152:641];
            r204 = r203[383:352];
            r205 = r202; r205[1024:993] = r204;
            // d.w[12] = q.w[12];
            //
            r206 = r1[1152:641];
            r207 = r206[415:384];
            r208 = r205; r208[1056:1025] = r207;
            // d.w[13] = q.w[13];
            //
            r209 = r1[1152:641];
            r210 = r209[447:416];
            r211 = r208; r211[1088:1057] = r210;
            // d.w[14] = q.w[14];
            //
            r212 = r1[1152:641];
            r213 = r212[479:448];
            r214 = r211; r214[1120:1089] = r213;
            // d.w[15] = q.w[15];
            //
            r215 = r1[1152:641];
            r216 = r215[511:480];
            r217 = r214; r217[1152:1121] = r216;
            r218 = (r60) ? (r169) : (r217);
            // if round_val < 64 {
            //    let current_w = if round_val < 16 {
            //       let idx = round_val as b64;
            //       if idx == 0 {
            //          q.w[0]
            //       }
            //        else if idx == 1 {
            //          q.w[1]
            //       }
            //        else if idx == 2 {
            //          q.w[2]
            //       }
            //        else if idx == 3 {
            //          q.w[3]
            //       }
            //        else if idx == 4 {
            //          q.w[4]
            //       }
            //        else if idx == 5 {
            //          q.w[5]
            //       }
            //        else if idx == 6 {
            //          q.w[6]
            //       }
            //        else if idx == 7 {
            //          q.w[7]
            //       }
            //        else if idx == 8 {
            //          q.w[8]
            //       }
            //        else if idx == 9 {
            //          q.w[9]
            //       }
            //        else if idx == 10 {
            //          q.w[10]
            //       }
            //        else if idx == 11 {
            //          q.w[11]
            //       }
            //        else if idx == 12 {
            //          q.w[12]
            //       }
            //        else if idx == 13 {
            //          q.w[13]
            //       }
            //        else if idx == 14 {
            //          q.w[14]
            //       }
            //        else {
            //          q.w[15]
            //       }
            //
            //    }
            //     else {
            //       d.w[15]
            //    }
            //    ;
            //    let s1 = sigma1(q.state.e);
            //    let ch_result = ch(q.state.e, q.state.f, q.state.g);
            //    let temp1 = q.state.h_reg + s1 + ch_result + get_k(q.state.round) + current_w;
            //    let s0 = sigma0(q.state.a);
            //    let maj_result = maj(q.state.a, q.state.b, q.state.c);
            //    let temp2 = s0 + maj_result;
            //    d.state.h_reg = q.state.g;
            //    d.state.g = q.state.f;
            //    d.state.f = q.state.e;
            //    d.state.e = q.state.d + temp1;
            //    d.state.d = q.state.c;
            //    d.state.c = q.state.b;
            //    d.state.b = q.state.a;
            //    d.state.a = temp1 + temp2;
            //    d.state.round = bits(round_val + 1);
            //    if round_val == 63 {
            //       d.state.h[0] = q.state.h[0] + d.state.a;
            //       d.state.h[1] = q.state.h[1] + d.state.b;
            //       d.state.h[2] = q.state.h[2] + d.state.c;
            //       d.state.h[3] = q.state.h[3] + d.state.d;
            //       d.state.h[4] = q.state.h[4] + d.state.e;
            //       d.state.h[5] = q.state.h[5] + d.state.f;
            //       d.state.h[6] = q.state.h[6] + d.state.g;
            //       d.state.h[7] = q.state.h[7] + d.state.h_reg;
            //       d.state.done = true;
            //       output_valid = true;
            //       hash_out = d.state.h;
            //    }
            //
            // }
            //
            //
            r219 = r57 < l18;
            // let current_w = if round_val < 16 {
            //    let idx = round_val as b64;
            //    if idx == 0 {
            //       q.w[0]
            //    }
            //     else if idx == 1 {
            //       q.w[1]
            //    }
            //     else if idx == 2 {
            //       q.w[2]
            //    }
            //     else if idx == 3 {
            //       q.w[3]
            //    }
            //     else if idx == 4 {
            //       q.w[4]
            //    }
            //     else if idx == 5 {
            //       q.w[5]
            //    }
            //     else if idx == 6 {
            //       q.w[6]
            //    }
            //     else if idx == 7 {
            //       q.w[7]
            //    }
            //     else if idx == 8 {
            //       q.w[8]
            //    }
            //     else if idx == 9 {
            //       q.w[9]
            //    }
            //     else if idx == 10 {
            //       q.w[10]
            //    }
            //     else if idx == 11 {
            //       q.w[11]
            //    }
            //     else if idx == 12 {
            //       q.w[12]
            //    }
            //     else if idx == 13 {
            //       q.w[13]
            //    }
            //     else if idx == 14 {
            //       q.w[14]
            //    }
            //     else {
            //       q.w[15]
            //    }
            //
            // }
            //  else {
            //    d.w[15]
            // }
            // ;
            //
            r220 = r57 < l19;
            // let idx = round_val as b64;
            //
            r221 = r57[63:0];
            // if idx == 0 {
            //    q.w[0]
            // }
            //  else if idx == 1 {
            //    q.w[1]
            // }
            //  else if idx == 2 {
            //    q.w[2]
            // }
            //  else if idx == 3 {
            //    q.w[3]
            // }
            //  else if idx == 4 {
            //    q.w[4]
            // }
            //  else if idx == 5 {
            //    q.w[5]
            // }
            //  else if idx == 6 {
            //    q.w[6]
            // }
            //  else if idx == 7 {
            //    q.w[7]
            // }
            //  else if idx == 8 {
            //    q.w[8]
            // }
            //  else if idx == 9 {
            //    q.w[9]
            // }
            //  else if idx == 10 {
            //    q.w[10]
            // }
            //  else if idx == 11 {
            //    q.w[11]
            // }
            //  else if idx == 12 {
            //    q.w[12]
            // }
            //  else if idx == 13 {
            //    q.w[13]
            // }
            //  else if idx == 14 {
            //    q.w[14]
            // }
            //  else {
            //    q.w[15]
            // }
            //
            //
            r222 = r221 == l20;
            // q.w[0]
            //
            r223 = r1[1152:641];
            r224 = r223[31:0];
            r225 = r221 == l21;
            // q.w[1]
            //
            r226 = r1[1152:641];
            r227 = r226[63:32];
            r228 = r221 == l22;
            // q.w[2]
            //
            r229 = r1[1152:641];
            r230 = r229[95:64];
            r231 = r221 == l23;
            // q.w[3]
            //
            r232 = r1[1152:641];
            r233 = r232[127:96];
            r234 = r221 == l24;
            // q.w[4]
            //
            r235 = r1[1152:641];
            r236 = r235[159:128];
            r237 = r221 == l25;
            // q.w[5]
            //
            r238 = r1[1152:641];
            r239 = r238[191:160];
            r240 = r221 == l26;
            // q.w[6]
            //
            r241 = r1[1152:641];
            r242 = r241[223:192];
            r243 = r221 == l27;
            // q.w[7]
            //
            r244 = r1[1152:641];
            r245 = r244[255:224];
            r246 = r221 == l28;
            // q.w[8]
            //
            r247 = r1[1152:641];
            r248 = r247[287:256];
            r249 = r221 == l29;
            // q.w[9]
            //
            r250 = r1[1152:641];
            r251 = r250[319:288];
            r252 = r221 == l30;
            // q.w[10]
            //
            r253 = r1[1152:641];
            r254 = r253[351:320];
            r255 = r221 == l31;
            // q.w[11]
            //
            r256 = r1[1152:641];
            r257 = r256[383:352];
            r258 = r221 == l32;
            // q.w[12]
            //
            r259 = r1[1152:641];
            r260 = r259[415:384];
            r261 = r221 == l33;
            // q.w[13]
            //
            r262 = r1[1152:641];
            r263 = r262[447:416];
            r264 = r221 == l34;
            // q.w[14]
            //
            r265 = r1[1152:641];
            r266 = r265[479:448];
            // q.w[15]
            //
            r267 = r1[1152:641];
            r268 = r267[511:480];
            r269 = (r264) ? (r266) : (r268);
            r270 = (r261) ? (r263) : (r269);
            r271 = (r258) ? (r260) : (r270);
            r272 = (r255) ? (r257) : (r271);
            r273 = (r252) ? (r254) : (r272);
            r274 = (r249) ? (r251) : (r273);
            r275 = (r246) ? (r248) : (r274);
            r276 = (r243) ? (r245) : (r275);
            r277 = (r240) ? (r242) : (r276);
            r278 = (r237) ? (r239) : (r277);
            r279 = (r234) ? (r236) : (r278);
            r280 = (r231) ? (r233) : (r279);
            r281 = (r228) ? (r230) : (r280);
            r282 = (r225) ? (r227) : (r281);
            r283 = (r222) ? (r224) : (r282);
            // d.w[15]
            //
            r284 = r218[1152:641];
            r285 = r284[511:480];
            r286 = (r220) ? (r283) : (r285);
            // let s1 = sigma1(q.state.e);
            //
            r287 = r1[640:0];
            r288 = r287[415:384];
            // rotr(x, 6) ^ rotr(x, 11) ^ rotr(x, 25)
            //
            // let n = n & 31;
            //
            // (x >> n) | (x << (32 - n))
            //
            r558 = { {6{1'b0}}, r288 };
            r294 = r558[37:6];
            r568 = r288[5:0];
            r296 = { r568, l90 };
            r297 = r294 | r296;
            // let n = n & 31;
            //
            // (x >> n) | (x << (32 - n))
            //
            r559 = { {11{1'b0}}, r288 };
            r302 = r559[42:11];
            r569 = r288[10:0];
            r304 = { r569, l91 };
            r305 = r302 | r304;
            r307 = r297 ^ r305;
            // let n = n & 31;
            //
            // (x >> n) | (x << (32 - n))
            //
            r560 = { {25{1'b0}}, r288 };
            r311 = r560[56:25];
            r570 = r288[24:0];
            r313 = { r570, l92 };
            r314 = r311 | r313;
            r290 = r307 ^ r314;
            // let ch_result = ch(q.state.e, q.state.f, q.state.g);
            //
            r317 = r1[640:0];
            r318 = r317[415:384];
            r319 = r1[640:0];
            r320 = r319[447:416];
            r321 = r1[640:0];
            r322 = r321[479:448];
            // (x & y) ^ (!x & z)
            //
            r327 = r318 & r320;
            r328 = ~(r318);
            r329 = r328 & r322;
            r326 = r327 ^ r329;
            // let temp1 = q.state.h_reg + s1 + ch_result + get_k(q.state.round) + current_w;
            //
            r331 = r1[640:0];
            r332 = r331[511:480];
            r333 = r332 + r290;
            r334 = r333 + r326;
            r335 = r1[640:0];
            r336 = r335[639:512];
            // let r = round.raw() as b64;
            //
            r339 = r336[63:0];
            // if r < 64 {
            //    bits(K[r])
            // }
            //  else {
            //    bits(0)
            // }
            //
            //
            r340 = r339 < l44;
            // bits(K[r])
            //
            r341 = r339[13:0];
            r550 = { {14{1'b0}}, r341 };
            r553 = r550[20:0];
            r342 = { r553, l65 };
            r343 = r342[13:0];
            r344 = l46 + r343;
            r345 = l47[(r344) +: 128];
            r346 = r345[31:0];
            // bits(0)
            //
            r338 = (r340) ? (r346) : (l48);
            r348 = r334 + r338;
            r349 = r348 + r286;
            // let s0 = sigma0(q.state.a);
            //
            r350 = r1[640:0];
            r351 = r350[287:256];
            // rotr(x, 2) ^ rotr(x, 13) ^ rotr(x, 22)
            //
            // let n = n & 31;
            //
            // (x >> n) | (x << (32 - n))
            //
            r561 = { {2{1'b0}}, r351 };
            r357 = r561[33:2];
            r571 = r351[1:0];
            r359 = { r571, l93 };
            r360 = r357 | r359;
            // let n = n & 31;
            //
            // (x >> n) | (x << (32 - n))
            //
            r562 = { {13{1'b0}}, r351 };
            r365 = r562[44:13];
            r572 = r351[12:0];
            r367 = { r572, l94 };
            r368 = r365 | r367;
            r370 = r360 ^ r368;
            // let n = n & 31;
            //
            // (x >> n) | (x << (32 - n))
            //
            r563 = { {22{1'b0}}, r351 };
            r374 = r563[53:22];
            r573 = r351[21:0];
            r376 = { r573, l95 };
            r377 = r374 | r376;
            r353 = r370 ^ r377;
            // let maj_result = maj(q.state.a, q.state.b, q.state.c);
            //
            r380 = r1[640:0];
            r381 = r380[287:256];
            r382 = r1[640:0];
            r383 = r382[319:288];
            r384 = r1[640:0];
            r385 = r384[351:320];
            // (x & y) ^ (x & z) ^ (y & z)
            //
            r390 = r381 & r383;
            r391 = r381 & r385;
            r392 = r390 ^ r391;
            r393 = r383 & r385;
            r389 = r392 ^ r393;
            // let temp2 = s0 + maj_result;
            //
            r395 = r353 + r389;
            // d.state.h_reg = q.state.g;
            //
            r396 = r1[640:0];
            r397 = r396[479:448];
            r398 = r218; r398[511:480] = r397;
            // d.state.g = q.state.f;
            //
            r399 = r1[640:0];
            r400 = r399[447:416];
            r401 = r398; r401[479:448] = r400;
            // d.state.f = q.state.e;
            //
            r402 = r1[640:0];
            r403 = r402[415:384];
            r404 = r401; r404[447:416] = r403;
            // d.state.e = q.state.d + temp1;
            //
            r405 = r1[640:0];
            r406 = r405[383:352];
            r407 = r406 + r349;
            r408 = r404; r408[415:384] = r407;
            // d.state.d = q.state.c;
            //
            r409 = r1[640:0];
            r410 = r409[351:320];
            r411 = r408; r411[383:352] = r410;
            // d.state.c = q.state.b;
            //
            r412 = r1[640:0];
            r413 = r412[319:288];
            r414 = r411; r414[351:320] = r413;
            // d.state.b = q.state.a;
            //
            r415 = r1[640:0];
            r416 = r415[287:256];
            r417 = r414; r417[319:288] = r416;
            // d.state.a = temp1 + temp2;
            //
            r418 = r349 + r395;
            r419 = r417; r419[287:256] = r418;
            // d.state.round = bits(round_val + 1);
            //
            r420 = r57 + l58;
            r421 = r420[127:0];
            r422 = r419; r422[639:512] = r421;
            // if round_val == 63 {
            //    d.state.h[0] = q.state.h[0] + d.state.a;
            //    d.state.h[1] = q.state.h[1] + d.state.b;
            //    d.state.h[2] = q.state.h[2] + d.state.c;
            //    d.state.h[3] = q.state.h[3] + d.state.d;
            //    d.state.h[4] = q.state.h[4] + d.state.e;
            //    d.state.h[5] = q.state.h[5] + d.state.f;
            //    d.state.h[6] = q.state.h[6] + d.state.g;
            //    d.state.h[7] = q.state.h[7] + d.state.h_reg;
            //    d.state.done = true;
            //    output_valid = true;
            //    hash_out = d.state.h;
            // }
            //
            //
            r423 = r57 == l59;
            // d.state.h[0] = q.state.h[0] + d.state.a;
            //
            r424 = r1[640:0];
            r425 = r424[255:0];
            r426 = r425[31:0];
            r427 = r422[640:0];
            r428 = r427[287:256];
            r429 = r426 + r428;
            r430 = r422; r430[31:0] = r429;
            // d.state.h[1] = q.state.h[1] + d.state.b;
            //
            r431 = r1[640:0];
            r432 = r431[255:0];
            r433 = r432[63:32];
            r434 = r430[640:0];
            r435 = r434[319:288];
            r436 = r433 + r435;
            r437 = r430; r437[63:32] = r436;
            // d.state.h[2] = q.state.h[2] + d.state.c;
            //
            r438 = r1[640:0];
            r439 = r438[255:0];
            r440 = r439[95:64];
            r441 = r437[640:0];
            r442 = r441[351:320];
            r443 = r440 + r442;
            r444 = r437; r444[95:64] = r443;
            // d.state.h[3] = q.state.h[3] + d.state.d;
            //
            r445 = r1[640:0];
            r446 = r445[255:0];
            r447 = r446[127:96];
            r448 = r444[640:0];
            r449 = r448[383:352];
            r450 = r447 + r449;
            r451 = r444; r451[127:96] = r450;
            // d.state.h[4] = q.state.h[4] + d.state.e;
            //
            r452 = r1[640:0];
            r453 = r452[255:0];
            r454 = r453[159:128];
            r455 = r451[640:0];
            r456 = r455[415:384];
            r457 = r454 + r456;
            r458 = r451; r458[159:128] = r457;
            // d.state.h[5] = q.state.h[5] + d.state.f;
            //
            r459 = r1[640:0];
            r460 = r459[255:0];
            r461 = r460[191:160];
            r462 = r458[640:0];
            r463 = r462[447:416];
            r464 = r461 + r463;
            r465 = r458; r465[191:160] = r464;
            // d.state.h[6] = q.state.h[6] + d.state.g;
            //
            r466 = r1[640:0];
            r467 = r466[255:0];
            r468 = r467[223:192];
            r469 = r465[640:0];
            r470 = r469[479:448];
            r471 = r468 + r470;
            r472 = r465; r472[223:192] = r471;
            // d.state.h[7] = q.state.h[7] + d.state.h_reg;
            //
            r473 = r1[640:0];
            r474 = r473[255:0];
            r475 = r474[255:224];
            r476 = r472[640:0];
            r477 = r476[511:480];
            r478 = r475 + r477;
            r479 = r472; r479[255:224] = r478;
            // d.state.done = true;
            //
            r480 = r479; r480[640:640] = l60;
            // output_valid = true;
            //
            // hash_out = d.state.h;
            //
            r481 = r480[640:0];
            r482 = r481[255:0];
            r483 = (r423) ? (r480) : (r422);
            r484 = (r423) ? (r482) : (r2);
            r485 = (r423) ? (l61) : (l62);
            r486 = (r219) ? (r483) : (r218);
            r487 = (r219) ? (r484) : (r2);
            r488 = (r219) ? (r485) : (l62);
            // d.state = q.state;
            //
            r489 = r1[640:0];
            r490 = l1; r490[640:0] = r489;
            // d.w[0] = q.w[0];
            //
            r491 = r1[1152:641];
            r492 = r491[31:0];
            r493 = r490; r493[672:641] = r492;
            // d.w[1] = q.w[1];
            //
            r494 = r1[1152:641];
            r495 = r494[63:32];
            r496 = r493; r496[704:673] = r495;
            // d.w[2] = q.w[2];
            //
            r497 = r1[1152:641];
            r498 = r497[95:64];
            r499 = r496; r499[736:705] = r498;
            // d.w[3] = q.w[3];
            //
            r500 = r1[1152:641];
            r501 = r500[127:96];
            r502 = r499; r502[768:737] = r501;
            // d.w[4] = q.w[4];
            //
            r503 = r1[1152:641];
            r504 = r503[159:128];
            r505 = r502; r505[800:769] = r504;
            // d.w[5] = q.w[5];
            //
            r506 = r1[1152:641];
            r507 = r506[191:160];
            r508 = r505; r508[832:801] = r507;
            // d.w[6] = q.w[6];
            //
            r509 = r1[1152:641];
            r510 = r509[223:192];
            r511 = r508; r511[864:833] = r510;
            // d.w[7] = q.w[7];
            //
            r512 = r1[1152:641];
            r513 = r512[255:224];
            r514 = r511; r514[896:865] = r513;
            // d.w[8] = q.w[8];
            //
            r515 = r1[1152:641];
            r516 = r515[287:256];
            r517 = r514; r517[928:897] = r516;
            // d.w[9] = q.w[9];
            //
            r518 = r1[1152:641];
            r519 = r518[319:288];
            r520 = r517; r520[960:929] = r519;
            // d.w[10] = q.w[10];
            //
            r521 = r1[1152:641];
            r522 = r521[351:320];
            r523 = r520; r523[992:961] = r522;
            // d.w[11] = q.w[11];
            //
            r524 = r1[1152:641];
            r525 = r524[383:352];
            r526 = r523; r526[1024:993] = r525;
            // d.w[12] = q.w[12];
            //
            r527 = r1[1152:641];
            r528 = r527[415:384];
            r529 = r526; r529[1056:1025] = r528;
            // d.w[13] = q.w[13];
            //
            r530 = r1[1152:641];
            r531 = r530[447:416];
            r532 = r529; r532[1088:1057] = r531;
            // d.w[14] = q.w[14];
            //
            r533 = r1[1152:641];
            r534 = r533[479:448];
            r535 = r532; r535[1120:1089] = r534;
            // d.w[15] = q.w[15];
            //
            r536 = r1[1152:641];
            r537 = r536[511:480];
            r538 = r535; r538[1152:1121] = r537;
            // output_valid = true;
            //
            // hash_out = q.state.h;
            //
            r539 = r1[640:0];
            r540 = r539[255:0];
            r541 = (r55) ? (r486) : (r538);
            r542 = (r55) ? (r487) : (r540);
            r543 = (r55) ? (r488) : (l63);
            r544 = (r3) ? (r52) : (r541);
            r545 = (r3) ? (r2) : (r542);
            r546 = (r3) ? (l62) : (r543);
            // ((hash_out, output_valid, ), d, )
            //
            r547 = { r546, r545 };
            r548 = { r544, r547 };
            kernel_kernel = r548;
        end
    endfunction
endmodule
//
module top_state(input wire [1:0] clock_reset, input wire [640:0] i, output reg [640:0] o);
    wire [0:0] clock;
    wire [0:0] reset;
    initial begin
        o = 641'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    assign clock = clock_reset[0];
    assign reset = clock_reset[1];
    always @(posedge clock) begin
        if (reset)
        begin
            o <= 641'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        end else begin
            o <= i;
        end
    end
endmodule
// array of 16 x Positive edge triggered DFF holding value of type b32, with reset value of 0_b32
module top_w(input wire [1:0] clock_reset, input wire [511:0] i, output wire [511:0] o);
    top_w_0 c0 (.clock_reset(clock_reset),.i(i[31:0]),.o(o[31:0]));
    top_w_1 c1 (.clock_reset(clock_reset),.i(i[63:32]),.o(o[63:32]));
    top_w_10 c2 (.clock_reset(clock_reset),.i(i[95:64]),.o(o[95:64]));
    top_w_11 c3 (.clock_reset(clock_reset),.i(i[127:96]),.o(o[127:96]));
    top_w_12 c4 (.clock_reset(clock_reset),.i(i[159:128]),.o(o[159:128]));
    top_w_13 c5 (.clock_reset(clock_reset),.i(i[191:160]),.o(o[191:160]));
    top_w_14 c6 (.clock_reset(clock_reset),.i(i[223:192]),.o(o[223:192]));
    top_w_15 c7 (.clock_reset(clock_reset),.i(i[255:224]),.o(o[255:224]));
    top_w_2 c8 (.clock_reset(clock_reset),.i(i[287:256]),.o(o[287:256]));
    top_w_3 c9 (.clock_reset(clock_reset),.i(i[319:288]),.o(o[319:288]));
    top_w_4 c10 (.clock_reset(clock_reset),.i(i[351:320]),.o(o[351:320]));
    top_w_5 c11 (.clock_reset(clock_reset),.i(i[383:352]),.o(o[383:352]));
    top_w_6 c12 (.clock_reset(clock_reset),.i(i[415:384]),.o(o[415:384]));
    top_w_7 c13 (.clock_reset(clock_reset),.i(i[447:416]),.o(o[447:416]));
    top_w_8 c14 (.clock_reset(clock_reset),.i(i[479:448]),.o(o[479:448]));
    top_w_9 c15 (.clock_reset(clock_reset),.i(i[511:480]),.o(o[511:480]));
endmodule
//
module top_w_0(input wire [1:0] clock_reset, input wire [31:0] i, output reg [31:0] o);
    wire [0:0] clock;
    wire [0:0] reset;
    initial begin
        o = 32'b00000000000000000000000000000000;
    end
    assign clock = clock_reset[0];
    assign reset = clock_reset[1];
    always @(posedge clock) begin
        if (reset)
        begin
            o <= 32'b00000000000000000000000000000000;
        end else begin
            o <= i;
        end
    end
endmodule
//
module top_w_1(input wire [1:0] clock_reset, input wire [31:0] i, output reg [31:0] o);
    wire [0:0] clock;
    wire [0:0] reset;
    initial begin
        o = 32'b00000000000000000000000000000000;
    end
    assign clock = clock_reset[0];
    assign reset = clock_reset[1];
    always @(posedge clock) begin
        if (reset)
        begin
            o <= 32'b00000000000000000000000000000000;
        end else begin
            o <= i;
        end
    end
endmodule
//
module top_w_10(input wire [1:0] clock_reset, input wire [31:0] i, output reg [31:0] o);
    wire [0:0] clock;
    wire [0:0] reset;
    initial begin
        o = 32'b00000000000000000000000000000000;
    end
    assign clock = clock_reset[0];
    assign reset = clock_reset[1];
    always @(posedge clock) begin
        if (reset)
        begin
            o <= 32'b00000000000000000000000000000000;
        end else begin
            o <= i;
        end
    end
endmodule
//
module top_w_11(input wire [1:0] clock_reset, input wire [31:0] i, output reg [31:0] o);
    wire [0:0] clock;
    wire [0:0] reset;
    initial begin
        o = 32'b00000000000000000000000000000000;
    end
    assign clock = clock_reset[0];
    assign reset = clock_reset[1];
    always @(posedge clock) begin
        if (reset)
        begin
            o <= 32'b00000000000000000000000000000000;
        end else begin
            o <= i;
        end
    end
endmodule
//
module top_w_12(input wire [1:0] clock_reset, input wire [31:0] i, output reg [31:0] o);
    wire [0:0] clock;
    wire [0:0] reset;
    initial begin
        o = 32'b00000000000000000000000000000000;
    end
    assign clock = clock_reset[0];
    assign reset = clock_reset[1];
    always @(posedge clock) begin
        if (reset)
        begin
            o <= 32'b00000000000000000000000000000000;
        end else begin
            o <= i;
        end
    end
endmodule
//
module top_w_13(input wire [1:0] clock_reset, input wire [31:0] i, output reg [31:0] o);
    wire [0:0] clock;
    wire [0:0] reset;
    initial begin
        o = 32'b00000000000000000000000000000000;
    end
    assign clock = clock_reset[0];
    assign reset = clock_reset[1];
    always @(posedge clock) begin
        if (reset)
        begin
            o <= 32'b00000000000000000000000000000000;
        end else begin
            o <= i;
        end
    end
endmodule
//
module top_w_14(input wire [1:0] clock_reset, input wire [31:0] i, output reg [31:0] o);
    wire [0:0] clock;
    wire [0:0] reset;
    initial begin
        o = 32'b00000000000000000000000000000000;
    end
    assign clock = clock_reset[0];
    assign reset = clock_reset[1];
    always @(posedge clock) begin
        if (reset)
        begin
            o <= 32'b00000000000000000000000000000000;
        end else begin
            o <= i;
        end
    end
endmodule
//
module top_w_15(input wire [1:0] clock_reset, input wire [31:0] i, output reg [31:0] o);
    wire [0:0] clock;
    wire [0:0] reset;
    initial begin
        o = 32'b00000000000000000000000000000000;
    end
    assign clock = clock_reset[0];
    assign reset = clock_reset[1];
    always @(posedge clock) begin
        if (reset)
        begin
            o <= 32'b00000000000000000000000000000000;
        end else begin
            o <= i;
        end
    end
endmodule
//
module top_w_2(input wire [1:0] clock_reset, input wire [31:0] i, output reg [31:0] o);
    wire [0:0] clock;
    wire [0:0] reset;
    initial begin
        o = 32'b00000000000000000000000000000000;
    end
    assign clock = clock_reset[0];
    assign reset = clock_reset[1];
    always @(posedge clock) begin
        if (reset)
        begin
            o <= 32'b00000000000000000000000000000000;
        end else begin
            o <= i;
        end
    end
endmodule
//
module top_w_3(input wire [1:0] clock_reset, input wire [31:0] i, output reg [31:0] o);
    wire [0:0] clock;
    wire [0:0] reset;
    initial begin
        o = 32'b00000000000000000000000000000000;
    end
    assign clock = clock_reset[0];
    assign reset = clock_reset[1];
    always @(posedge clock) begin
        if (reset)
        begin
            o <= 32'b00000000000000000000000000000000;
        end else begin
            o <= i;
        end
    end
endmodule
//
module top_w_4(input wire [1:0] clock_reset, input wire [31:0] i, output reg [31:0] o);
    wire [0:0] clock;
    wire [0:0] reset;
    initial begin
        o = 32'b00000000000000000000000000000000;
    end
    assign clock = clock_reset[0];
    assign reset = clock_reset[1];
    always @(posedge clock) begin
        if (reset)
        begin
            o <= 32'b00000000000000000000000000000000;
        end else begin
            o <= i;
        end
    end
endmodule
//
module top_w_5(input wire [1:0] clock_reset, input wire [31:0] i, output reg [31:0] o);
    wire [0:0] clock;
    wire [0:0] reset;
    initial begin
        o = 32'b00000000000000000000000000000000;
    end
    assign clock = clock_reset[0];
    assign reset = clock_reset[1];
    always @(posedge clock) begin
        if (reset)
        begin
            o <= 32'b00000000000000000000000000000000;
        end else begin
            o <= i;
        end
    end
endmodule
//
module top_w_6(input wire [1:0] clock_reset, input wire [31:0] i, output reg [31:0] o);
    wire [0:0] clock;
    wire [0:0] reset;
    initial begin
        o = 32'b00000000000000000000000000000000;
    end
    assign clock = clock_reset[0];
    assign reset = clock_reset[1];
    always @(posedge clock) begin
        if (reset)
        begin
            o <= 32'b00000000000000000000000000000000;
        end else begin
            o <= i;
        end
    end
endmodule
//
module top_w_7(input wire [1:0] clock_reset, input wire [31:0] i, output reg [31:0] o);
    wire [0:0] clock;
    wire [0:0] reset;
    initial begin
        o = 32'b00000000000000000000000000000000;
    end
    assign clock = clock_reset[0];
    assign reset = clock_reset[1];
    always @(posedge clock) begin
        if (reset)
        begin
            o <= 32'b00000000000000000000000000000000;
        end else begin
            o <= i;
        end
    end
endmodule
//
module top_w_8(input wire [1:0] clock_reset, input wire [31:0] i, output reg [31:0] o);
    wire [0:0] clock;
    wire [0:0] reset;
    initial begin
        o = 32'b00000000000000000000000000000000;
    end
    assign clock = clock_reset[0];
    assign reset = clock_reset[1];
    always @(posedge clock) begin
        if (reset)
        begin
            o <= 32'b00000000000000000000000000000000;
        end else begin
            o <= i;
        end
    end
endmodule
//
module top_w_9(input wire [1:0] clock_reset, input wire [31:0] i, output reg [31:0] o);
    wire [0:0] clock;
    wire [0:0] reset;
    initial begin
        o = 32'b00000000000000000000000000000000;
    end
    assign clock = clock_reset[0];
    assign reset = clock_reset[1];
    always @(posedge clock) begin
        if (reset)
        begin
            o <= 32'b00000000000000000000000000000000;
        end else begin
            o <= i;
        end
    end
endmodule
